
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"dc",x"fb",x"c2",x"78"),
     1 => (x"c8",x"78",x"c0",x"48"),
     2 => (x"87",x"c5",x"02",x"66"),
     3 => (x"c2",x"49",x"ff",x"c3"),
     4 => (x"c2",x"49",x"c0",x"87"),
     5 => (x"cc",x"59",x"e4",x"fb"),
     6 => (x"87",x"c6",x"02",x"66"),
     7 => (x"4a",x"d5",x"d5",x"c5"),
     8 => (x"ff",x"cf",x"87",x"c4"),
     9 => (x"fb",x"c2",x"4a",x"ff"),
    10 => (x"fb",x"c2",x"5a",x"e8"),
    11 => (x"78",x"c1",x"48",x"e8"),
    12 => (x"4f",x"26",x"4b",x"26"),
    13 => (x"5c",x"5b",x"5e",x"0e"),
    14 => (x"4d",x"71",x"0e",x"5d"),
    15 => (x"bf",x"e4",x"fb",x"c2"),
    16 => (x"02",x"9d",x"75",x"4b"),
    17 => (x"c8",x"49",x"87",x"cb"),
    18 => (x"dc",x"ff",x"c1",x"91"),
    19 => (x"c4",x"82",x"71",x"4a"),
    20 => (x"dc",x"c3",x"c2",x"87"),
    21 => (x"12",x"4c",x"c0",x"4a"),
    22 => (x"c2",x"99",x"73",x"49"),
    23 => (x"48",x"bf",x"e0",x"fb"),
    24 => (x"d4",x"ff",x"b8",x"71"),
    25 => (x"b7",x"c1",x"78",x"08"),
    26 => (x"b7",x"c8",x"84",x"2b"),
    27 => (x"87",x"e7",x"04",x"ac"),
    28 => (x"bf",x"dc",x"fb",x"c2"),
    29 => (x"c2",x"80",x"c8",x"48"),
    30 => (x"26",x"58",x"e0",x"fb"),
    31 => (x"26",x"4c",x"26",x"4d"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"4b",x"71",x"1e",x"73"),
    34 => (x"02",x"9a",x"4a",x"13"),
    35 => (x"49",x"72",x"87",x"cb"),
    36 => (x"13",x"87",x"e1",x"fe"),
    37 => (x"f5",x"05",x"9a",x"4a"),
    38 => (x"26",x"4b",x"26",x"87"),
    39 => (x"fb",x"c2",x"1e",x"4f"),
    40 => (x"c2",x"49",x"bf",x"dc"),
    41 => (x"c1",x"48",x"dc",x"fb"),
    42 => (x"c0",x"c4",x"78",x"a1"),
    43 => (x"db",x"03",x"a9",x"b7"),
    44 => (x"48",x"d4",x"ff",x"87"),
    45 => (x"bf",x"e0",x"fb",x"c2"),
    46 => (x"dc",x"fb",x"c2",x"78"),
    47 => (x"fb",x"c2",x"49",x"bf"),
    48 => (x"a1",x"c1",x"48",x"dc"),
    49 => (x"b7",x"c0",x"c4",x"78"),
    50 => (x"87",x"e5",x"04",x"a9"),
    51 => (x"c8",x"48",x"d0",x"ff"),
    52 => (x"e8",x"fb",x"c2",x"78"),
    53 => (x"26",x"78",x"c0",x"48"),
    54 => (x"00",x"00",x"00",x"4f"),
    55 => (x"00",x"00",x"00",x"00"),
    56 => (x"00",x"00",x"00",x"00"),
    57 => (x"5f",x"00",x"00",x"00"),
    58 => (x"00",x"00",x"00",x"5f"),
    59 => (x"00",x"03",x"03",x"00"),
    60 => (x"00",x"00",x"03",x"03"),
    61 => (x"14",x"7f",x"7f",x"14"),
    62 => (x"00",x"14",x"7f",x"7f"),
    63 => (x"6b",x"2e",x"24",x"00"),
    64 => (x"00",x"12",x"3a",x"6b"),
    65 => (x"18",x"36",x"6a",x"4c"),
    66 => (x"00",x"32",x"56",x"6c"),
    67 => (x"59",x"4f",x"7e",x"30"),
    68 => (x"40",x"68",x"3a",x"77"),
    69 => (x"07",x"04",x"00",x"00"),
    70 => (x"00",x"00",x"00",x"03"),
    71 => (x"3e",x"1c",x"00",x"00"),
    72 => (x"00",x"00",x"41",x"63"),
    73 => (x"63",x"41",x"00",x"00"),
    74 => (x"00",x"00",x"1c",x"3e"),
    75 => (x"1c",x"3e",x"2a",x"08"),
    76 => (x"08",x"2a",x"3e",x"1c"),
    77 => (x"3e",x"08",x"08",x"00"),
    78 => (x"00",x"08",x"08",x"3e"),
    79 => (x"e0",x"80",x"00",x"00"),
    80 => (x"00",x"00",x"00",x"60"),
    81 => (x"08",x"08",x"08",x"00"),
    82 => (x"00",x"08",x"08",x"08"),
    83 => (x"60",x"00",x"00",x"00"),
    84 => (x"00",x"00",x"00",x"60"),
    85 => (x"18",x"30",x"60",x"40"),
    86 => (x"01",x"03",x"06",x"0c"),
    87 => (x"59",x"7f",x"3e",x"00"),
    88 => (x"00",x"3e",x"7f",x"4d"),
    89 => (x"7f",x"06",x"04",x"00"),
    90 => (x"00",x"00",x"00",x"7f"),
    91 => (x"71",x"63",x"42",x"00"),
    92 => (x"00",x"46",x"4f",x"59"),
    93 => (x"49",x"63",x"22",x"00"),
    94 => (x"00",x"36",x"7f",x"49"),
    95 => (x"13",x"16",x"1c",x"18"),
    96 => (x"00",x"10",x"7f",x"7f"),
    97 => (x"45",x"67",x"27",x"00"),
    98 => (x"00",x"39",x"7d",x"45"),
    99 => (x"4b",x"7e",x"3c",x"00"),
   100 => (x"00",x"30",x"79",x"49"),
   101 => (x"71",x"01",x"01",x"00"),
   102 => (x"00",x"07",x"0f",x"79"),
   103 => (x"49",x"7f",x"36",x"00"),
   104 => (x"00",x"36",x"7f",x"49"),
   105 => (x"49",x"4f",x"06",x"00"),
   106 => (x"00",x"1e",x"3f",x"69"),
   107 => (x"66",x"00",x"00",x"00"),
   108 => (x"00",x"00",x"00",x"66"),
   109 => (x"e6",x"80",x"00",x"00"),
   110 => (x"00",x"00",x"00",x"66"),
   111 => (x"14",x"08",x"08",x"00"),
   112 => (x"00",x"22",x"22",x"14"),
   113 => (x"14",x"14",x"14",x"00"),
   114 => (x"00",x"14",x"14",x"14"),
   115 => (x"14",x"22",x"22",x"00"),
   116 => (x"00",x"08",x"08",x"14"),
   117 => (x"51",x"03",x"02",x"00"),
   118 => (x"00",x"06",x"0f",x"59"),
   119 => (x"5d",x"41",x"7f",x"3e"),
   120 => (x"00",x"1e",x"1f",x"55"),
   121 => (x"09",x"7f",x"7e",x"00"),
   122 => (x"00",x"7e",x"7f",x"09"),
   123 => (x"49",x"7f",x"7f",x"00"),
   124 => (x"00",x"36",x"7f",x"49"),
   125 => (x"63",x"3e",x"1c",x"00"),
   126 => (x"00",x"41",x"41",x"41"),
   127 => (x"41",x"7f",x"7f",x"00"),
   128 => (x"00",x"1c",x"3e",x"63"),
   129 => (x"49",x"7f",x"7f",x"00"),
   130 => (x"00",x"41",x"41",x"49"),
   131 => (x"09",x"7f",x"7f",x"00"),
   132 => (x"00",x"01",x"01",x"09"),
   133 => (x"41",x"7f",x"3e",x"00"),
   134 => (x"00",x"7a",x"7b",x"49"),
   135 => (x"08",x"7f",x"7f",x"00"),
   136 => (x"00",x"7f",x"7f",x"08"),
   137 => (x"7f",x"41",x"00",x"00"),
   138 => (x"00",x"00",x"41",x"7f"),
   139 => (x"40",x"60",x"20",x"00"),
   140 => (x"00",x"3f",x"7f",x"40"),
   141 => (x"1c",x"08",x"7f",x"7f"),
   142 => (x"00",x"41",x"63",x"36"),
   143 => (x"40",x"7f",x"7f",x"00"),
   144 => (x"00",x"40",x"40",x"40"),
   145 => (x"0c",x"06",x"7f",x"7f"),
   146 => (x"00",x"7f",x"7f",x"06"),
   147 => (x"0c",x"06",x"7f",x"7f"),
   148 => (x"00",x"7f",x"7f",x"18"),
   149 => (x"41",x"7f",x"3e",x"00"),
   150 => (x"00",x"3e",x"7f",x"41"),
   151 => (x"09",x"7f",x"7f",x"00"),
   152 => (x"00",x"06",x"0f",x"09"),
   153 => (x"61",x"41",x"7f",x"3e"),
   154 => (x"00",x"40",x"7e",x"7f"),
   155 => (x"09",x"7f",x"7f",x"00"),
   156 => (x"00",x"66",x"7f",x"19"),
   157 => (x"4d",x"6f",x"26",x"00"),
   158 => (x"00",x"32",x"7b",x"59"),
   159 => (x"7f",x"01",x"01",x"00"),
   160 => (x"00",x"01",x"01",x"7f"),
   161 => (x"40",x"7f",x"3f",x"00"),
   162 => (x"00",x"3f",x"7f",x"40"),
   163 => (x"70",x"3f",x"0f",x"00"),
   164 => (x"00",x"0f",x"3f",x"70"),
   165 => (x"18",x"30",x"7f",x"7f"),
   166 => (x"00",x"7f",x"7f",x"30"),
   167 => (x"1c",x"36",x"63",x"41"),
   168 => (x"41",x"63",x"36",x"1c"),
   169 => (x"7c",x"06",x"03",x"01"),
   170 => (x"01",x"03",x"06",x"7c"),
   171 => (x"4d",x"59",x"71",x"61"),
   172 => (x"00",x"41",x"43",x"47"),
   173 => (x"7f",x"7f",x"00",x"00"),
   174 => (x"00",x"00",x"41",x"41"),
   175 => (x"0c",x"06",x"03",x"01"),
   176 => (x"40",x"60",x"30",x"18"),
   177 => (x"41",x"41",x"00",x"00"),
   178 => (x"00",x"00",x"7f",x"7f"),
   179 => (x"03",x"06",x"0c",x"08"),
   180 => (x"00",x"08",x"0c",x"06"),
   181 => (x"80",x"80",x"80",x"80"),
   182 => (x"00",x"80",x"80",x"80"),
   183 => (x"03",x"00",x"00",x"00"),
   184 => (x"00",x"00",x"04",x"07"),
   185 => (x"54",x"74",x"20",x"00"),
   186 => (x"00",x"78",x"7c",x"54"),
   187 => (x"44",x"7f",x"7f",x"00"),
   188 => (x"00",x"38",x"7c",x"44"),
   189 => (x"44",x"7c",x"38",x"00"),
   190 => (x"00",x"00",x"44",x"44"),
   191 => (x"44",x"7c",x"38",x"00"),
   192 => (x"00",x"7f",x"7f",x"44"),
   193 => (x"54",x"7c",x"38",x"00"),
   194 => (x"00",x"18",x"5c",x"54"),
   195 => (x"7f",x"7e",x"04",x"00"),
   196 => (x"00",x"00",x"05",x"05"),
   197 => (x"a4",x"bc",x"18",x"00"),
   198 => (x"00",x"7c",x"fc",x"a4"),
   199 => (x"04",x"7f",x"7f",x"00"),
   200 => (x"00",x"78",x"7c",x"04"),
   201 => (x"3d",x"00",x"00",x"00"),
   202 => (x"00",x"00",x"40",x"7d"),
   203 => (x"80",x"80",x"80",x"00"),
   204 => (x"00",x"00",x"7d",x"fd"),
   205 => (x"10",x"7f",x"7f",x"00"),
   206 => (x"00",x"44",x"6c",x"38"),
   207 => (x"3f",x"00",x"00",x"00"),
   208 => (x"00",x"00",x"40",x"7f"),
   209 => (x"18",x"0c",x"7c",x"7c"),
   210 => (x"00",x"78",x"7c",x"0c"),
   211 => (x"04",x"7c",x"7c",x"00"),
   212 => (x"00",x"78",x"7c",x"04"),
   213 => (x"44",x"7c",x"38",x"00"),
   214 => (x"00",x"38",x"7c",x"44"),
   215 => (x"24",x"fc",x"fc",x"00"),
   216 => (x"00",x"18",x"3c",x"24"),
   217 => (x"24",x"3c",x"18",x"00"),
   218 => (x"00",x"fc",x"fc",x"24"),
   219 => (x"04",x"7c",x"7c",x"00"),
   220 => (x"00",x"08",x"0c",x"04"),
   221 => (x"54",x"5c",x"48",x"00"),
   222 => (x"00",x"20",x"74",x"54"),
   223 => (x"7f",x"3f",x"04",x"00"),
   224 => (x"00",x"00",x"44",x"44"),
   225 => (x"40",x"7c",x"3c",x"00"),
   226 => (x"00",x"7c",x"7c",x"40"),
   227 => (x"60",x"3c",x"1c",x"00"),
   228 => (x"00",x"1c",x"3c",x"60"),
   229 => (x"30",x"60",x"7c",x"3c"),
   230 => (x"00",x"3c",x"7c",x"60"),
   231 => (x"10",x"38",x"6c",x"44"),
   232 => (x"00",x"44",x"6c",x"38"),
   233 => (x"e0",x"bc",x"1c",x"00"),
   234 => (x"00",x"1c",x"3c",x"60"),
   235 => (x"74",x"64",x"44",x"00"),
   236 => (x"00",x"44",x"4c",x"5c"),
   237 => (x"3e",x"08",x"08",x"00"),
   238 => (x"00",x"41",x"41",x"77"),
   239 => (x"7f",x"00",x"00",x"00"),
   240 => (x"00",x"00",x"00",x"7f"),
   241 => (x"77",x"41",x"41",x"00"),
   242 => (x"00",x"08",x"08",x"3e"),
   243 => (x"03",x"01",x"01",x"02"),
   244 => (x"00",x"01",x"02",x"02"),
   245 => (x"7f",x"7f",x"7f",x"7f"),
   246 => (x"00",x"7f",x"7f",x"7f"),
   247 => (x"1c",x"1c",x"08",x"08"),
   248 => (x"7f",x"7f",x"3e",x"3e"),
   249 => (x"3e",x"3e",x"7f",x"7f"),
   250 => (x"08",x"08",x"1c",x"1c"),
   251 => (x"7c",x"18",x"10",x"00"),
   252 => (x"00",x"10",x"18",x"7c"),
   253 => (x"7c",x"30",x"10",x"00"),
   254 => (x"00",x"10",x"30",x"7c"),
   255 => (x"60",x"60",x"30",x"10"),
   256 => (x"00",x"06",x"1e",x"78"),
   257 => (x"18",x"3c",x"66",x"42"),
   258 => (x"00",x"42",x"66",x"3c"),
   259 => (x"c2",x"6a",x"38",x"78"),
   260 => (x"00",x"38",x"6c",x"c6"),
   261 => (x"60",x"00",x"00",x"60"),
   262 => (x"00",x"60",x"00",x"00"),
   263 => (x"5c",x"5b",x"5e",x"0e"),
   264 => (x"86",x"fc",x"0e",x"5d"),
   265 => (x"c2",x"59",x"a6",x"c4"),
   266 => (x"4c",x"bf",x"f0",x"fb"),
   267 => (x"1e",x"c0",x"4b",x"c0"),
   268 => (x"02",x"ab",x"66",x"c4"),
   269 => (x"4d",x"c0",x"87",x"c4"),
   270 => (x"4d",x"c1",x"87",x"c2"),
   271 => (x"49",x"73",x"1e",x"75"),
   272 => (x"c8",x"87",x"e0",x"ee"),
   273 => (x"49",x"e0",x"c0",x"86"),
   274 => (x"c4",x"87",x"e9",x"ef"),
   275 => (x"49",x"6a",x"4a",x"a4"),
   276 => (x"f1",x"87",x"f0",x"f0"),
   277 => (x"84",x"cc",x"87",x"c7"),
   278 => (x"b7",x"c8",x"83",x"c1"),
   279 => (x"cd",x"ff",x"04",x"ab"),
   280 => (x"26",x"8e",x"fc",x"87"),
   281 => (x"26",x"4c",x"26",x"4d"),
   282 => (x"1e",x"4f",x"26",x"4b"),
   283 => (x"fb",x"c2",x"4a",x"71"),
   284 => (x"fb",x"c2",x"5a",x"f4"),
   285 => (x"78",x"c7",x"48",x"f4"),
   286 => (x"87",x"e0",x"fe",x"49"),
   287 => (x"73",x"1e",x"4f",x"26"),
   288 => (x"fc",x"4b",x"71",x"1e"),
   289 => (x"73",x"0b",x"7b",x"0b"),
   290 => (x"c1",x"9a",x"c1",x"4a"),
   291 => (x"ed",x"49",x"a2",x"c0"),
   292 => (x"df",x"c2",x"87",x"c4"),
   293 => (x"4b",x"26",x"5b",x"f4"),
   294 => (x"71",x"1e",x"4f",x"26"),
   295 => (x"1e",x"66",x"c4",x"4a"),
   296 => (x"ca",x"ec",x"49",x"72"),
   297 => (x"26",x"8e",x"fc",x"87"),
   298 => (x"d4",x"ff",x"1e",x"4f"),
   299 => (x"78",x"ff",x"c3",x"48"),
   300 => (x"c0",x"48",x"d0",x"ff"),
   301 => (x"d4",x"ff",x"78",x"e1"),
   302 => (x"71",x"78",x"c1",x"48"),
   303 => (x"ff",x"30",x"c4",x"48"),
   304 => (x"ff",x"78",x"08",x"d4"),
   305 => (x"e0",x"c0",x"48",x"d0"),
   306 => (x"0e",x"4f",x"26",x"78"),
   307 => (x"5d",x"5c",x"5b",x"5e"),
   308 => (x"c8",x"86",x"ec",x"0e"),
   309 => (x"78",x"c0",x"48",x"a6"),
   310 => (x"bf",x"ec",x"80",x"c4"),
   311 => (x"c2",x"80",x"f8",x"78"),
   312 => (x"78",x"bf",x"f0",x"fb"),
   313 => (x"bf",x"f8",x"fb",x"c2"),
   314 => (x"4d",x"bf",x"e8",x"4c"),
   315 => (x"bf",x"f0",x"df",x"c2"),
   316 => (x"87",x"c1",x"e4",x"49"),
   317 => (x"fe",x"e8",x"49",x"c7"),
   318 => (x"c2",x"49",x"70",x"87"),
   319 => (x"87",x"d0",x"05",x"99"),
   320 => (x"bf",x"e8",x"df",x"c2"),
   321 => (x"cc",x"b9",x"ff",x"49"),
   322 => (x"99",x"c1",x"99",x"66"),
   323 => (x"87",x"cd",x"c2",x"02"),
   324 => (x"ff",x"48",x"a6",x"c8"),
   325 => (x"c7",x"78",x"bf",x"c8"),
   326 => (x"87",x"db",x"e8",x"49"),
   327 => (x"a6",x"c4",x"49",x"70"),
   328 => (x"05",x"99",x"71",x"5c"),
   329 => (x"66",x"cc",x"87",x"ce"),
   330 => (x"c4",x"99",x"c1",x"49"),
   331 => (x"99",x"71",x"5c",x"a6"),
   332 => (x"87",x"c4",x"c1",x"02"),
   333 => (x"c8",x"4c",x"c8",x"ff"),
   334 => (x"a6",x"cc",x"4b",x"66"),
   335 => (x"78",x"bf",x"ec",x"48"),
   336 => (x"cc",x"87",x"f2",x"e2"),
   337 => (x"48",x"6c",x"5b",x"a6"),
   338 => (x"a6",x"d4",x"88",x"73"),
   339 => (x"a8",x"e8",x"cf",x"58"),
   340 => (x"c2",x"87",x"d1",x"06"),
   341 => (x"49",x"bf",x"e4",x"df"),
   342 => (x"df",x"c2",x"b9",x"c1"),
   343 => (x"fd",x"71",x"59",x"e8"),
   344 => (x"4b",x"6c",x"87",x"c7"),
   345 => (x"ce",x"e7",x"49",x"c7"),
   346 => (x"05",x"98",x"70",x"87"),
   347 => (x"cc",x"87",x"cb",x"ff"),
   348 => (x"99",x"c1",x"49",x"66"),
   349 => (x"87",x"c2",x"ff",x"05"),
   350 => (x"df",x"c2",x"4c",x"6e"),
   351 => (x"c1",x"4a",x"bf",x"f0"),
   352 => (x"f4",x"df",x"c2",x"ba"),
   353 => (x"7a",x"0a",x"fc",x"5a"),
   354 => (x"c1",x"9a",x"c1",x"0a"),
   355 => (x"e9",x"49",x"a2",x"c0"),
   356 => (x"da",x"c1",x"87",x"c4"),
   357 => (x"87",x"df",x"e6",x"49"),
   358 => (x"c1",x"48",x"a6",x"c8"),
   359 => (x"e8",x"df",x"c2",x"78"),
   360 => (x"78",x"66",x"cc",x"48"),
   361 => (x"bf",x"f0",x"df",x"c2"),
   362 => (x"87",x"c7",x"c1",x"05"),
   363 => (x"4b",x"c0",x"c0",x"c8"),
   364 => (x"7e",x"d4",x"df",x"c2"),
   365 => (x"49",x"14",x"4c",x"6e"),
   366 => (x"70",x"87",x"fc",x"e5"),
   367 => (x"c2",x"c0",x"02",x"98"),
   368 => (x"c1",x"b5",x"73",x"87"),
   369 => (x"ff",x"05",x"2b",x"b7"),
   370 => (x"49",x"75",x"87",x"ec"),
   371 => (x"71",x"99",x"ff",x"c3"),
   372 => (x"fb",x"49",x"c0",x"1e"),
   373 => (x"49",x"75",x"87",x"c4"),
   374 => (x"71",x"29",x"b7",x"c8"),
   375 => (x"fa",x"49",x"c1",x"1e"),
   376 => (x"86",x"c8",x"87",x"f8"),
   377 => (x"e5",x"49",x"fd",x"c3"),
   378 => (x"fa",x"c3",x"87",x"cd"),
   379 => (x"87",x"c7",x"e5",x"49"),
   380 => (x"75",x"87",x"d2",x"c7"),
   381 => (x"99",x"ff",x"c3",x"49"),
   382 => (x"71",x"2d",x"b7",x"c8"),
   383 => (x"02",x"9d",x"75",x"b5"),
   384 => (x"ff",x"87",x"e0",x"c0"),
   385 => (x"6e",x"7e",x"bf",x"c8"),
   386 => (x"ec",x"df",x"c2",x"49"),
   387 => (x"e0",x"c2",x"89",x"bf"),
   388 => (x"c5",x"c0",x"03",x"a9"),
   389 => (x"c0",x"4d",x"c0",x"87"),
   390 => (x"df",x"c2",x"87",x"cf"),
   391 => (x"78",x"6e",x"48",x"ec"),
   392 => (x"c2",x"87",x"c6",x"c0"),
   393 => (x"c0",x"48",x"ec",x"df"),
   394 => (x"c8",x"49",x"75",x"78"),
   395 => (x"ce",x"c0",x"05",x"99"),
   396 => (x"49",x"f5",x"c3",x"87"),
   397 => (x"70",x"87",x"c0",x"e4"),
   398 => (x"02",x"99",x"c2",x"49"),
   399 => (x"c2",x"87",x"eb",x"c0"),
   400 => (x"02",x"bf",x"f4",x"fb"),
   401 => (x"48",x"87",x"ca",x"c0"),
   402 => (x"fb",x"c2",x"88",x"c1"),
   403 => (x"d4",x"c0",x"58",x"f8"),
   404 => (x"48",x"66",x"c4",x"87"),
   405 => (x"c4",x"80",x"e0",x"c1"),
   406 => (x"bf",x"6e",x"58",x"a6"),
   407 => (x"87",x"c5",x"c0",x"02"),
   408 => (x"73",x"49",x"ff",x"4b"),
   409 => (x"48",x"a6",x"c8",x"0f"),
   410 => (x"49",x"75",x"78",x"c1"),
   411 => (x"c0",x"05",x"99",x"c4"),
   412 => (x"f2",x"c3",x"87",x"ce"),
   413 => (x"87",x"ff",x"e2",x"49"),
   414 => (x"99",x"c2",x"49",x"70"),
   415 => (x"87",x"f2",x"c0",x"02"),
   416 => (x"bf",x"f4",x"fb",x"c2"),
   417 => (x"c7",x"48",x"6e",x"7e"),
   418 => (x"c0",x"03",x"a8",x"b7"),
   419 => (x"48",x"6e",x"87",x"cb"),
   420 => (x"fb",x"c2",x"80",x"c1"),
   421 => (x"d4",x"c0",x"58",x"f8"),
   422 => (x"48",x"66",x"c4",x"87"),
   423 => (x"c4",x"80",x"e0",x"c1"),
   424 => (x"bf",x"6e",x"58",x"a6"),
   425 => (x"87",x"c5",x"c0",x"02"),
   426 => (x"73",x"49",x"fe",x"4b"),
   427 => (x"48",x"a6",x"c8",x"0f"),
   428 => (x"fd",x"c3",x"78",x"c1"),
   429 => (x"87",x"ff",x"e1",x"49"),
   430 => (x"99",x"c2",x"49",x"70"),
   431 => (x"87",x"e6",x"c0",x"02"),
   432 => (x"bf",x"f4",x"fb",x"c2"),
   433 => (x"87",x"c9",x"c0",x"02"),
   434 => (x"48",x"f4",x"fb",x"c2"),
   435 => (x"d0",x"c0",x"78",x"c0"),
   436 => (x"4a",x"66",x"c4",x"87"),
   437 => (x"6a",x"82",x"e0",x"c1"),
   438 => (x"87",x"c5",x"c0",x"02"),
   439 => (x"73",x"49",x"fd",x"4b"),
   440 => (x"48",x"a6",x"c8",x"0f"),
   441 => (x"fa",x"c3",x"78",x"c1"),
   442 => (x"87",x"cb",x"e1",x"49"),
   443 => (x"99",x"c2",x"49",x"70"),
   444 => (x"87",x"ee",x"c0",x"02"),
   445 => (x"bf",x"f4",x"fb",x"c2"),
   446 => (x"a8",x"b7",x"c7",x"48"),
   447 => (x"87",x"c9",x"c0",x"03"),
   448 => (x"48",x"f4",x"fb",x"c2"),
   449 => (x"d4",x"c0",x"78",x"c7"),
   450 => (x"48",x"66",x"c4",x"87"),
   451 => (x"c4",x"80",x"e0",x"c1"),
   452 => (x"bf",x"6e",x"58",x"a6"),
   453 => (x"87",x"c5",x"c0",x"02"),
   454 => (x"73",x"49",x"fc",x"4b"),
   455 => (x"48",x"a6",x"c8",x"0f"),
   456 => (x"48",x"75",x"78",x"c1"),
   457 => (x"c4",x"98",x"f0",x"c3"),
   458 => (x"98",x"70",x"58",x"a6"),
   459 => (x"87",x"ce",x"c0",x"05"),
   460 => (x"e0",x"49",x"da",x"c1"),
   461 => (x"49",x"70",x"87",x"c1"),
   462 => (x"c1",x"02",x"99",x"c2"),
   463 => (x"05",x"6e",x"87",x"ca"),
   464 => (x"c1",x"87",x"cd",x"c0"),
   465 => (x"df",x"ff",x"49",x"da"),
   466 => (x"98",x"70",x"87",x"ed"),
   467 => (x"87",x"e8",x"c0",x"02"),
   468 => (x"4b",x"49",x"bf",x"e8"),
   469 => (x"c8",x"9b",x"ff",x"c3"),
   470 => (x"b3",x"71",x"29",x"b7"),
   471 => (x"87",x"d5",x"da",x"ff"),
   472 => (x"f0",x"c3",x"49",x"73"),
   473 => (x"05",x"99",x"71",x"99"),
   474 => (x"c1",x"87",x"e5",x"ff"),
   475 => (x"df",x"ff",x"49",x"da"),
   476 => (x"98",x"70",x"87",x"c5"),
   477 => (x"87",x"d8",x"ff",x"05"),
   478 => (x"bf",x"f4",x"fb",x"c2"),
   479 => (x"93",x"cc",x"4b",x"49"),
   480 => (x"6b",x"83",x"66",x"c4"),
   481 => (x"0f",x"73",x"71",x"4b"),
   482 => (x"c0",x"02",x"9c",x"74"),
   483 => (x"02",x"6c",x"87",x"e9"),
   484 => (x"6c",x"87",x"e4",x"c0"),
   485 => (x"de",x"de",x"ff",x"49"),
   486 => (x"c1",x"49",x"70",x"87"),
   487 => (x"cb",x"c0",x"02",x"99"),
   488 => (x"4b",x"a4",x"c4",x"87"),
   489 => (x"bf",x"f4",x"fb",x"c2"),
   490 => (x"0f",x"4b",x"6b",x"49"),
   491 => (x"c0",x"02",x"84",x"c8"),
   492 => (x"05",x"6c",x"87",x"c5"),
   493 => (x"c8",x"87",x"dc",x"ff"),
   494 => (x"c8",x"c0",x"02",x"66"),
   495 => (x"f4",x"fb",x"c2",x"87"),
   496 => (x"d7",x"f1",x"49",x"bf"),
   497 => (x"26",x"8e",x"ec",x"87"),
   498 => (x"26",x"4c",x"26",x"4d"),
   499 => (x"00",x"4f",x"26",x"4b"),
   500 => (x"00",x"00",x"00",x"10"),
   501 => (x"14",x"11",x"12",x"58"),
   502 => (x"23",x"1c",x"1b",x"1d"),
   503 => (x"94",x"91",x"59",x"5a"),
   504 => (x"f4",x"eb",x"f2",x"f5"),
   505 => (x"00",x"00",x"00",x"00"),
   506 => (x"00",x"00",x"00",x"00"),
   507 => (x"00",x"00",x"00",x"00"),
   508 => (x"00",x"00",x"00",x"00"),
   509 => (x"5c",x"5b",x"5e",x"0e"),
   510 => (x"4b",x"71",x"0e",x"5d"),
   511 => (x"d0",x"4c",x"d4",x"ff"),
   512 => (x"78",x"c0",x"48",x"66"),
   513 => (x"dd",x"ff",x"49",x"d6"),
   514 => (x"ff",x"c3",x"87",x"ea"),
   515 => (x"c3",x"49",x"6c",x"7c"),
   516 => (x"4d",x"71",x"99",x"ff"),
   517 => (x"99",x"f0",x"c3",x"49"),
   518 => (x"05",x"a9",x"e0",x"c1"),
   519 => (x"ff",x"c3",x"87",x"cb"),
   520 => (x"c3",x"48",x"6c",x"7c"),
   521 => (x"08",x"66",x"d0",x"98"),
   522 => (x"7c",x"ff",x"c3",x"78"),
   523 => (x"c8",x"49",x"4a",x"6c"),
   524 => (x"7c",x"ff",x"c3",x"31"),
   525 => (x"b2",x"71",x"4a",x"6c"),
   526 => (x"31",x"c8",x"49",x"72"),
   527 => (x"6c",x"7c",x"ff",x"c3"),
   528 => (x"72",x"b2",x"71",x"4a"),
   529 => (x"c3",x"31",x"c8",x"49"),
   530 => (x"4a",x"6c",x"7c",x"ff"),
   531 => (x"d0",x"ff",x"b2",x"71"),
   532 => (x"78",x"e0",x"c0",x"48"),
   533 => (x"c2",x"02",x"9b",x"73"),
   534 => (x"75",x"7b",x"72",x"87"),
   535 => (x"26",x"4d",x"26",x"48"),
   536 => (x"26",x"4b",x"26",x"4c"),
   537 => (x"4f",x"26",x"1e",x"4f"),
   538 => (x"5c",x"5b",x"5e",x"0e"),
   539 => (x"76",x"86",x"f8",x"0e"),
   540 => (x"80",x"c4",x"48",x"1e"),
   541 => (x"fb",x"fd",x"49",x"70"),
   542 => (x"70",x"86",x"c4",x"87"),
   543 => (x"c3",x"48",x"6e",x"4b"),
   544 => (x"f4",x"c2",x"01",x"a8"),
   545 => (x"c3",x"4a",x"73",x"87"),
   546 => (x"d0",x"c1",x"9a",x"f0"),
   547 => (x"87",x"c7",x"02",x"aa"),
   548 => (x"05",x"aa",x"e0",x"c1"),
   549 => (x"73",x"87",x"e2",x"c2"),
   550 => (x"02",x"99",x"c8",x"49"),
   551 => (x"c4",x"ff",x"87",x"c3"),
   552 => (x"c3",x"4c",x"73",x"87"),
   553 => (x"05",x"ac",x"c2",x"9c"),
   554 => (x"c4",x"87",x"c4",x"c1"),
   555 => (x"31",x"c9",x"49",x"66"),
   556 => (x"66",x"c4",x"1e",x"71"),
   557 => (x"92",x"cc",x"c1",x"4a"),
   558 => (x"49",x"fc",x"fb",x"c2"),
   559 => (x"cc",x"fe",x"81",x"72"),
   560 => (x"49",x"d8",x"87",x"fa"),
   561 => (x"87",x"ec",x"da",x"ff"),
   562 => (x"c2",x"1e",x"c0",x"c8"),
   563 => (x"fd",x"49",x"f4",x"e8"),
   564 => (x"ff",x"87",x"cc",x"e6"),
   565 => (x"e0",x"c0",x"48",x"d0"),
   566 => (x"f4",x"e8",x"c2",x"78"),
   567 => (x"4a",x"66",x"cc",x"1e"),
   568 => (x"c2",x"92",x"cc",x"c1"),
   569 => (x"72",x"49",x"fc",x"fb"),
   570 => (x"d0",x"cb",x"fe",x"81"),
   571 => (x"c1",x"86",x"cc",x"87"),
   572 => (x"c4",x"c1",x"05",x"ac"),
   573 => (x"49",x"66",x"c4",x"87"),
   574 => (x"1e",x"71",x"31",x"c9"),
   575 => (x"c1",x"4a",x"66",x"c4"),
   576 => (x"fb",x"c2",x"92",x"cc"),
   577 => (x"81",x"72",x"49",x"fc"),
   578 => (x"87",x"f0",x"cb",x"fe"),
   579 => (x"1e",x"f4",x"e8",x"c2"),
   580 => (x"c1",x"4a",x"66",x"c8"),
   581 => (x"fb",x"c2",x"92",x"cc"),
   582 => (x"81",x"72",x"49",x"fc"),
   583 => (x"87",x"de",x"c9",x"fe"),
   584 => (x"d9",x"ff",x"49",x"d7"),
   585 => (x"c0",x"c8",x"87",x"ce"),
   586 => (x"f4",x"e8",x"c2",x"1e"),
   587 => (x"cb",x"e4",x"fd",x"49"),
   588 => (x"ff",x"86",x"cc",x"87"),
   589 => (x"e0",x"c0",x"48",x"d0"),
   590 => (x"26",x"8e",x"f8",x"78"),
   591 => (x"26",x"4b",x"26",x"4c"),
   592 => (x"4a",x"71",x"1e",x"4f"),
   593 => (x"03",x"aa",x"b7",x"c4"),
   594 => (x"49",x"72",x"87",x"ce"),
   595 => (x"c2",x"91",x"cc",x"c1"),
   596 => (x"c1",x"81",x"fc",x"fb"),
   597 => (x"79",x"c0",x"81",x"c8"),
   598 => (x"5e",x"0e",x"4f",x"26"),
   599 => (x"0e",x"5d",x"5c",x"5b"),
   600 => (x"4a",x"71",x"86",x"fc"),
   601 => (x"c0",x"4b",x"d4",x"ff"),
   602 => (x"4d",x"66",x"d4",x"4c"),
   603 => (x"01",x"ad",x"b7",x"c3"),
   604 => (x"72",x"87",x"c2",x"c2"),
   605 => (x"ec",x"c0",x"02",x"9a"),
   606 => (x"49",x"75",x"1e",x"87"),
   607 => (x"c2",x"91",x"cc",x"c1"),
   608 => (x"71",x"48",x"fc",x"fb"),
   609 => (x"58",x"a6",x"c8",x"80"),
   610 => (x"fe",x"49",x"66",x"c4"),
   611 => (x"c4",x"87",x"f9",x"c2"),
   612 => (x"02",x"98",x"70",x"86"),
   613 => (x"49",x"6e",x"87",x"d4"),
   614 => (x"c1",x"81",x"c8",x"c1"),
   615 => (x"c8",x"49",x"6e",x"79"),
   616 => (x"c5",x"4c",x"69",x"81"),
   617 => (x"fe",x"49",x"75",x"87"),
   618 => (x"d0",x"ff",x"87",x"d7"),
   619 => (x"78",x"e1",x"c8",x"48"),
   620 => (x"48",x"74",x"7b",x"dd"),
   621 => (x"70",x"98",x"ff",x"c3"),
   622 => (x"c8",x"49",x"74",x"7b"),
   623 => (x"48",x"71",x"29",x"b7"),
   624 => (x"70",x"98",x"ff",x"c3"),
   625 => (x"d0",x"49",x"74",x"7b"),
   626 => (x"48",x"71",x"29",x"b7"),
   627 => (x"70",x"98",x"ff",x"c3"),
   628 => (x"d8",x"48",x"74",x"7b"),
   629 => (x"7b",x"70",x"28",x"b7"),
   630 => (x"7b",x"7b",x"7b",x"c0"),
   631 => (x"7b",x"7b",x"7b",x"7b"),
   632 => (x"7b",x"7b",x"7b",x"7b"),
   633 => (x"48",x"d0",x"ff",x"7b"),
   634 => (x"75",x"78",x"e0",x"c0"),
   635 => (x"ff",x"49",x"dc",x"1e"),
   636 => (x"c4",x"87",x"e6",x"d6"),
   637 => (x"26",x"8e",x"fc",x"86"),
   638 => (x"26",x"4c",x"26",x"4d"),
   639 => (x"14",x"4f",x"26",x"4b"),
   640 => (x"14",x"00",x"00",x"1d"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

