library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4c0c387",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49c4c0c3",
    18 => x"48dce7c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"d9e7c287",
    25 => x"d5e7c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"edc187f7",
    29 => x"e7c287fc",
    30 => x"e7c24dd9",
    31 => x"ad744cd9",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"5c5b5e0e",
    36 => x"86f00e5d",
    37 => x"a6c44cc0",
    38 => x"c078c048",
    39 => x"c04ba6e4",
    40 => x"484966e0",
    41 => x"e4c080c1",
    42 => x"7e1158a6",
    43 => x"f1c3026e",
    44 => x"0266c487",
    45 => x"c487c6c3",
    46 => x"78c048a6",
    47 => x"f0c04a6e",
    48 => x"dac2028a",
    49 => x"8af3c087",
    50 => x"87dbc202",
    51 => x"dc028ac1",
    52 => x"028ac887",
    53 => x"c487c8c2",
    54 => x"87d1028a",
    55 => x"c1028ac3",
    56 => x"8ac287eb",
    57 => x"c387c602",
    58 => x"c9c2058a",
    59 => x"7383c487",
    60 => x"6989c449",
    61 => x"c1026e7e",
    62 => x"a6c887c8",
    63 => x"c478c048",
    64 => x"cc78c080",
    65 => x"4a6e4d66",
    66 => x"cf2ab7dc",
    67 => x"c4486e9a",
    68 => x"727e7030",
    69 => x"87c5029a",
    70 => x"c148a6c8",
    71 => x"06aac978",
    72 => x"f7c087c5",
    73 => x"c087c382",
    74 => x"66c882f0",
    75 => x"7287c702",
    76 => x"87fac149",
    77 => x"85c184c1",
    78 => x"04adb7c8",
    79 => x"c187c7ff",
    80 => x"f0c087ce",
    81 => x"87e6c149",
    82 => x"c3c184c1",
    83 => x"7383c487",
    84 => x"6a8ac44a",
    85 => x"87f1c149",
    86 => x"4ca44970",
    87 => x"c487f1c0",
    88 => x"78c148a6",
    89 => x"c487e9c0",
    90 => x"c44a7383",
    91 => x"c0496a8a",
    92 => x"84c187fc",
    93 => x"496e87da",
    94 => x"d387f3c0",
    95 => x"c0486e87",
    96 => x"c705a8e5",
    97 => x"48a6c487",
    98 => x"87c478c1",
    99 => x"87de496e",
   100 => x"4966e0c0",
   101 => x"c080c148",
   102 => x"1158a6e4",
   103 => x"fc056e7e",
   104 => x"487487cf",
   105 => x"4d268ef0",
   106 => x"4b264c26",
   107 => x"fc1e4f26",
   108 => x"ff4a7186",
   109 => x"486949c0",
   110 => x"7098c0c4",
   111 => x"0298487e",
   112 => x"797287f4",
   113 => x"268efc48",
   114 => x"5b5e0e4f",
   115 => x"4b710e5c",
   116 => x"4a134cc0",
   117 => x"87cd029a",
   118 => x"d1ff4972",
   119 => x"1384c187",
   120 => x"f3059a4a",
   121 => x"26487487",
   122 => x"264b264c",
   123 => x"1e721e4f",
   124 => x"48121e73",
   125 => x"87ca0211",
   126 => x"98dfc34b",
   127 => x"0288739b",
   128 => x"4b2687f0",
   129 => x"4f264a26",
   130 => x"721e731e",
   131 => x"048bc11e",
   132 => x"481287ca",
   133 => x"87c40211",
   134 => x"87f10288",
   135 => x"4b264a26",
   136 => x"731e4f26",
   137 => x"a9738148",
   138 => x"1287c502",
   139 => x"87f60553",
   140 => x"731e4f26",
   141 => x"c84a711e",
   142 => x"c1494b66",
   143 => x"0299718b",
   144 => x"481287cf",
   145 => x"7808d4ff",
   146 => x"8bc14973",
   147 => x"f1059971",
   148 => x"264b2687",
   149 => x"5b5e0e4f",
   150 => x"4a710e5c",
   151 => x"cc4cd4ff",
   152 => x"c1494b66",
   153 => x"0299718b",
   154 => x"ffc387ce",
   155 => x"73526c7c",
   156 => x"718bc149",
   157 => x"87f20599",
   158 => x"4b264c26",
   159 => x"731e4f26",
   160 => x"4bd4ff1e",
   161 => x"6b7bffc3",
   162 => x"7bffc34a",
   163 => x"32c8496b",
   164 => x"ffc3b172",
   165 => x"c84a6b7b",
   166 => x"c3b27131",
   167 => x"496b7bff",
   168 => x"b17232c8",
   169 => x"4b264871",
   170 => x"5e0e4f26",
   171 => x"0e5d5c5b",
   172 => x"d4ff4d71",
   173 => x"c348754c",
   174 => x"7c7098ff",
   175 => x"bfdce7c2",
   176 => x"d087c805",
   177 => x"30c94866",
   178 => x"d058a6d4",
   179 => x"29d84966",
   180 => x"ffc34871",
   181 => x"d07c7098",
   182 => x"29d04966",
   183 => x"ffc34871",
   184 => x"d07c7098",
   185 => x"29c84966",
   186 => x"ffc34871",
   187 => x"d07c7098",
   188 => x"ffc34866",
   189 => x"757c7098",
   190 => x"7129d049",
   191 => x"98ffc348",
   192 => x"4b6c7c70",
   193 => x"4afff0c9",
   194 => x"05abffc3",
   195 => x"714987cf",
   196 => x"c14b6c7c",
   197 => x"87c5028a",
   198 => x"f202ab71",
   199 => x"26487387",
   200 => x"264c264d",
   201 => x"1e4f264b",
   202 => x"d4ff49c0",
   203 => x"78ffc348",
   204 => x"c8c381c1",
   205 => x"f104a9b7",
   206 => x"0e4f2687",
   207 => x"5d5c5b5e",
   208 => x"f0ffc00e",
   209 => x"c14df7c1",
   210 => x"c0c0c0c0",
   211 => x"d6ff4bc0",
   212 => x"dff8c487",
   213 => x"751ec04c",
   214 => x"87cefd49",
   215 => x"a8c186c4",
   216 => x"87e5c005",
   217 => x"c348d4ff",
   218 => x"1e7378ff",
   219 => x"c1f0e1c0",
   220 => x"f5fc49e9",
   221 => x"7086c487",
   222 => x"87ca0598",
   223 => x"c348d4ff",
   224 => x"48c178ff",
   225 => x"defe87cb",
   226 => x"058cc187",
   227 => x"c087c6ff",
   228 => x"264d2648",
   229 => x"264b264c",
   230 => x"5b5e0e4f",
   231 => x"ffc00e5c",
   232 => x"4cc1c1f0",
   233 => x"c348d4ff",
   234 => x"dccf78ff",
   235 => x"87d9f849",
   236 => x"1ec04bd3",
   237 => x"f1fb4974",
   238 => x"7086c487",
   239 => x"87ca0598",
   240 => x"c348d4ff",
   241 => x"48c178ff",
   242 => x"dafd87cb",
   243 => x"058bc187",
   244 => x"c087dfff",
   245 => x"264c2648",
   246 => x"004f264b",
   247 => x"00444d43",
   248 => x"43484453",
   249 => x"69616620",
   250 => x"000a216c",
   251 => x"52524549",
   252 => x"00000000",
   253 => x"00495053",
   254 => x"74697257",
   255 => x"61662065",
   256 => x"64656c69",
   257 => x"5e0e000a",
   258 => x"0e5d5c5b",
   259 => x"ff4dffc3",
   260 => x"d2fc4bd4",
   261 => x"1eeac687",
   262 => x"c1f0e1c0",
   263 => x"c9fa49c8",
   264 => x"c186c487",
   265 => x"87c802a8",
   266 => x"c087eefd",
   267 => x"87e8c148",
   268 => x"7087cbf9",
   269 => x"ffffcf49",
   270 => x"a9eac699",
   271 => x"fd87c802",
   272 => x"48c087d7",
   273 => x"7587d1c1",
   274 => x"4cf1c07b",
   275 => x"7087ecfb",
   276 => x"ecc00298",
   277 => x"c01ec087",
   278 => x"fac1f0ff",
   279 => x"87caf949",
   280 => x"987086c4",
   281 => x"7587da05",
   282 => x"75496b7b",
   283 => x"757b757b",
   284 => x"c17b757b",
   285 => x"c40299c0",
   286 => x"db48c187",
   287 => x"d748c087",
   288 => x"05acc287",
   289 => x"e0cf87ca",
   290 => x"87fdf449",
   291 => x"87c848c0",
   292 => x"fe058cc1",
   293 => x"48c087f6",
   294 => x"4c264d26",
   295 => x"4f264b26",
   296 => x"5c5b5e0e",
   297 => x"d0ff0e5d",
   298 => x"d0e5c04d",
   299 => x"c24cc0c1",
   300 => x"c148dce7",
   301 => x"49f4cf78",
   302 => x"c787cef4",
   303 => x"f97dc24b",
   304 => x"7dc387e5",
   305 => x"49741ec0",
   306 => x"c487dff7",
   307 => x"05a8c186",
   308 => x"c24b87c1",
   309 => x"87cb05ab",
   310 => x"f349eccf",
   311 => x"48c087eb",
   312 => x"c187f6c0",
   313 => x"d4ff058b",
   314 => x"87dafc87",
   315 => x"58e0e7c2",
   316 => x"cd059870",
   317 => x"c01ec187",
   318 => x"d0c1f0ff",
   319 => x"87eaf649",
   320 => x"d4ff86c4",
   321 => x"78ffc348",
   322 => x"c287eec4",
   323 => x"c258e4e7",
   324 => x"48d4ff7d",
   325 => x"c178ffc3",
   326 => x"264d2648",
   327 => x"264b264c",
   328 => x"5b5e0e4f",
   329 => x"710e5d5c",
   330 => x"4cffc34d",
   331 => x"744bd4ff",
   332 => x"48d0ff7b",
   333 => x"7478c3c4",
   334 => x"c01e757b",
   335 => x"d8c1f0ff",
   336 => x"87e6f549",
   337 => x"987086c4",
   338 => x"cf87cb02",
   339 => x"f8f149f8",
   340 => x"c048c187",
   341 => x"7b7487ee",
   342 => x"c87bfec3",
   343 => x"66d41ec0",
   344 => x"87cef349",
   345 => x"7b7486c4",
   346 => x"7b747b74",
   347 => x"4ae0dad8",
   348 => x"056b7b74",
   349 => x"8ac187c5",
   350 => x"7487f505",
   351 => x"48d0ff7b",
   352 => x"48c078c2",
   353 => x"4c264d26",
   354 => x"4f264b26",
   355 => x"5c5b5e0e",
   356 => x"86fc0e5d",
   357 => x"d4ff4b71",
   358 => x"c57ec04c",
   359 => x"4adfcdee",
   360 => x"6c7cffc3",
   361 => x"a8fec348",
   362 => x"87f8c005",
   363 => x"9b734d74",
   364 => x"d487cc02",
   365 => x"49731e66",
   366 => x"c487daf2",
   367 => x"ff87d486",
   368 => x"d1c448d0",
   369 => x"4a66d478",
   370 => x"c17dffc3",
   371 => x"87f8058a",
   372 => x"c35aa6d8",
   373 => x"737c7cff",
   374 => x"87c5059b",
   375 => x"d048d0ff",
   376 => x"7e4ac178",
   377 => x"fe058ac1",
   378 => x"486e87f6",
   379 => x"4d268efc",
   380 => x"4b264c26",
   381 => x"731e4f26",
   382 => x"c04a711e",
   383 => x"48d4ff4b",
   384 => x"ff78ffc3",
   385 => x"c3c448d0",
   386 => x"48d4ff78",
   387 => x"7278ffc3",
   388 => x"f0ffc01e",
   389 => x"f249d1c1",
   390 => x"86c487d0",
   391 => x"d2059870",
   392 => x"1ec0c887",
   393 => x"fd4966cc",
   394 => x"86c487e2",
   395 => x"d0ff4b70",
   396 => x"7378c248",
   397 => x"264b2648",
   398 => x"5b5e0e4f",
   399 => x"c00e5d5c",
   400 => x"f0ffc01e",
   401 => x"f149c9c1",
   402 => x"1ed287e0",
   403 => x"49ece7c2",
   404 => x"c887f9fc",
   405 => x"c14cc086",
   406 => x"acb7d284",
   407 => x"c287f804",
   408 => x"bf97ece7",
   409 => x"99c0c349",
   410 => x"05a9c0c1",
   411 => x"c287e7c0",
   412 => x"bf97f3e7",
   413 => x"c231d049",
   414 => x"bf97f4e7",
   415 => x"7232c84a",
   416 => x"f5e7c2b1",
   417 => x"b14abf97",
   418 => x"ffcf4c71",
   419 => x"c19cffff",
   420 => x"c134ca84",
   421 => x"e7c287e7",
   422 => x"49bf97f5",
   423 => x"99c631c1",
   424 => x"97f6e7c2",
   425 => x"b7c74abf",
   426 => x"c2b1722a",
   427 => x"bf97f1e7",
   428 => x"9dcf4d4a",
   429 => x"97f2e7c2",
   430 => x"9ac34abf",
   431 => x"e7c232ca",
   432 => x"4bbf97f3",
   433 => x"b27333c2",
   434 => x"97f4e7c2",
   435 => x"c0c34bbf",
   436 => x"2bb7c69b",
   437 => x"81c2b273",
   438 => x"307148c1",
   439 => x"48c14970",
   440 => x"4d703075",
   441 => x"84c14c72",
   442 => x"c0c89471",
   443 => x"cc06adb7",
   444 => x"b734c187",
   445 => x"b7c0c82d",
   446 => x"f4ff01ad",
   447 => x"26487487",
   448 => x"264c264d",
   449 => x"0e4f264b",
   450 => x"5d5c5b5e",
   451 => x"c286fc0e",
   452 => x"c048d4f0",
   453 => x"cce8c278",
   454 => x"fb49c01e",
   455 => x"86c487d8",
   456 => x"c5059870",
   457 => x"c948c087",
   458 => x"4dc087d5",
   459 => x"48d0f5c2",
   460 => x"e9c278c1",
   461 => x"e6c04ac2",
   462 => x"4bc849d8",
   463 => x"7087c9eb",
   464 => x"87c60598",
   465 => x"48d0f5c2",
   466 => x"e9c278c0",
   467 => x"e6c04ade",
   468 => x"4bc849e4",
   469 => x"7087f1ea",
   470 => x"87c60598",
   471 => x"48d0f5c2",
   472 => x"f5c278c0",
   473 => x"c002bfd0",
   474 => x"efc287fe",
   475 => x"c24dbfd2",
   476 => x"bf9fcaf0",
   477 => x"c5486e7e",
   478 => x"05a8ead6",
   479 => x"efc287c7",
   480 => x"ce4dbfd2",
   481 => x"ca486e87",
   482 => x"02a8d5e9",
   483 => x"48c087c5",
   484 => x"c287ecc7",
   485 => x"751ecce8",
   486 => x"87daf949",
   487 => x"987086c4",
   488 => x"c087c505",
   489 => x"87d7c748",
   490 => x"4adee9c2",
   491 => x"49f0e6c0",
   492 => x"d3e94bc8",
   493 => x"05987087",
   494 => x"c287c8c0",
   495 => x"c148d4f0",
   496 => x"c287d878",
   497 => x"c04ac2e9",
   498 => x"c849fce6",
   499 => x"87f8e84b",
   500 => x"c0029870",
   501 => x"48c087c5",
   502 => x"c287e4c6",
   503 => x"bf97caf0",
   504 => x"a9d5c149",
   505 => x"87cdc005",
   506 => x"97cbf0c2",
   507 => x"eac249bf",
   508 => x"c5c002a9",
   509 => x"c648c087",
   510 => x"e8c287c5",
   511 => x"7ebf97cc",
   512 => x"e9c3486e",
   513 => x"cec002a8",
   514 => x"c3486e87",
   515 => x"c002a8eb",
   516 => x"48c087c5",
   517 => x"c287e8c5",
   518 => x"bf97d7e8",
   519 => x"c0059949",
   520 => x"e8c287cc",
   521 => x"49bf97d8",
   522 => x"c002a9c2",
   523 => x"48c087c5",
   524 => x"c287ccc5",
   525 => x"bf97d9e8",
   526 => x"d0f0c248",
   527 => x"484c7058",
   528 => x"f0c288c1",
   529 => x"e8c258d4",
   530 => x"49bf97da",
   531 => x"e8c28175",
   532 => x"4abf97db",
   533 => x"a17232c8",
   534 => x"ecf4c27e",
   535 => x"c2786e48",
   536 => x"bf97dce8",
   537 => x"c4f5c248",
   538 => x"d4f0c258",
   539 => x"d3c202bf",
   540 => x"dee9c287",
   541 => x"cce6c04a",
   542 => x"e64bc849",
   543 => x"987087ca",
   544 => x"87c5c002",
   545 => x"f6c348c0",
   546 => x"ccf0c287",
   547 => x"f5c24cbf",
   548 => x"e8c25cc0",
   549 => x"49bf97f1",
   550 => x"e8c231c8",
   551 => x"4abf97f0",
   552 => x"e8c249a1",
   553 => x"4abf97f2",
   554 => x"a17232d0",
   555 => x"f3e8c249",
   556 => x"d84abf97",
   557 => x"49a17232",
   558 => x"59c8f5c2",
   559 => x"bfc0f5c2",
   560 => x"ecf4c291",
   561 => x"f4c281bf",
   562 => x"e8c259f4",
   563 => x"4abf97f9",
   564 => x"e8c232c8",
   565 => x"4bbf97f8",
   566 => x"e8c24aa2",
   567 => x"4bbf97fa",
   568 => x"a27333d0",
   569 => x"fbe8c24a",
   570 => x"cf4bbf97",
   571 => x"7333d89b",
   572 => x"f4c24aa2",
   573 => x"8ac25af8",
   574 => x"f4c29274",
   575 => x"a17248f8",
   576 => x"87c7c178",
   577 => x"97dee8c2",
   578 => x"31c849bf",
   579 => x"97dde8c2",
   580 => x"49a14abf",
   581 => x"ffc731c5",
   582 => x"c229c981",
   583 => x"c259c0f5",
   584 => x"bf97e3e8",
   585 => x"c232c84a",
   586 => x"bf97e2e8",
   587 => x"c24aa24b",
   588 => x"c25ac8f5",
   589 => x"92bfc0f5",
   590 => x"f4c2826e",
   591 => x"f4c25afc",
   592 => x"78c048f4",
   593 => x"48f0f4c2",
   594 => x"c278a172",
   595 => x"c248c8f5",
   596 => x"78bff4f4",
   597 => x"48ccf5c2",
   598 => x"bff8f4c2",
   599 => x"d4f0c278",
   600 => x"c9c002bf",
   601 => x"c4487487",
   602 => x"c07e7030",
   603 => x"f4c287c9",
   604 => x"c448bffc",
   605 => x"c27e7030",
   606 => x"6e48d8f0",
   607 => x"fc48c178",
   608 => x"264d268e",
   609 => x"264b264c",
   610 => x"0000004f",
   611 => x"33544146",
   612 => x"20202032",
   613 => x"00000000",
   614 => x"31544146",
   615 => x"20202036",
   616 => x"00000000",
   617 => x"33544146",
   618 => x"20202032",
   619 => x"00000000",
   620 => x"33544146",
   621 => x"20202032",
   622 => x"00000000",
   623 => x"31544146",
   624 => x"20202036",
   625 => x"5b5e0e00",
   626 => x"710e5d5c",
   627 => x"d4f0c24a",
   628 => x"87cb02bf",
   629 => x"2bc74b72",
   630 => x"ffc14d72",
   631 => x"7287c99d",
   632 => x"722bc84b",
   633 => x"9dffc34d",
   634 => x"bfecf4c2",
   635 => x"d0fec083",
   636 => x"d902abbf",
   637 => x"d4fec087",
   638 => x"cce8c25b",
   639 => x"ef49731e",
   640 => x"86c487f4",
   641 => x"c5059870",
   642 => x"c048c087",
   643 => x"f0c287e6",
   644 => x"d202bfd4",
   645 => x"c4497587",
   646 => x"cce8c291",
   647 => x"cf4c6981",
   648 => x"ffffffff",
   649 => x"7587cb9c",
   650 => x"c291c249",
   651 => x"9f81cce8",
   652 => x"48744c69",
   653 => x"4c264d26",
   654 => x"4f264b26",
   655 => x"5c5b5e0e",
   656 => x"86f40e5d",
   657 => x"c459a6c8",
   658 => x"80c84866",
   659 => x"486e7e70",
   660 => x"c11e78c0",
   661 => x"87fdcc49",
   662 => x"4c7086c4",
   663 => x"fcc0029c",
   664 => x"dcf0c287",
   665 => x"4966dc4a",
   666 => x"87c1deff",
   667 => x"c0029870",
   668 => x"4a7487eb",
   669 => x"cb4966dc",
   670 => x"cbdeff4b",
   671 => x"02987087",
   672 => x"1ec087db",
   673 => x"c4029c74",
   674 => x"c24dc087",
   675 => x"754dc187",
   676 => x"87c1cc49",
   677 => x"4c7086c4",
   678 => x"c4ff059c",
   679 => x"029c7487",
   680 => x"dc87f4c1",
   681 => x"486e49a4",
   682 => x"a4da7869",
   683 => x"4d66c449",
   684 => x"699f85c4",
   685 => x"d4f0c27d",
   686 => x"87d202bf",
   687 => x"9f49a4d4",
   688 => x"ffc04969",
   689 => x"487199ff",
   690 => x"7e7030d0",
   691 => x"7ec087c2",
   692 => x"6d48496e",
   693 => x"c47d7080",
   694 => x"78c04866",
   695 => x"cc4966c4",
   696 => x"c4796d81",
   697 => x"81d04966",
   698 => x"a6c879c0",
   699 => x"c878c048",
   700 => x"66c44c66",
   701 => x"7482d44a",
   702 => x"7291c849",
   703 => x"41c049a1",
   704 => x"84c1796d",
   705 => x"04acb7c6",
   706 => x"c487e7ff",
   707 => x"c4c14966",
   708 => x"c179c081",
   709 => x"c087c248",
   710 => x"268ef448",
   711 => x"264c264d",
   712 => x"0e4f264b",
   713 => x"5d5c5b5e",
   714 => x"d04c710e",
   715 => x"496c4d66",
   716 => x"c2b97585",
   717 => x"4abfd0f0",
   718 => x"9972baff",
   719 => x"c0029971",
   720 => x"a4c487e4",
   721 => x"f9496b4b",
   722 => x"7b7087fb",
   723 => x"bfccf0c2",
   724 => x"71816c49",
   725 => x"c2b9757c",
   726 => x"4abfd0f0",
   727 => x"9972baff",
   728 => x"ff059971",
   729 => x"7c7587dc",
   730 => x"4c264d26",
   731 => x"4f264b26",
   732 => x"711e731e",
   733 => x"f0f4c24b",
   734 => x"a3c449bf",
   735 => x"c24a6a4a",
   736 => x"ccf0c28a",
   737 => x"a17292bf",
   738 => x"d0f0c249",
   739 => x"9a6b4abf",
   740 => x"c049a172",
   741 => x"c859d4fe",
   742 => x"e9711e66",
   743 => x"86c487d8",
   744 => x"c4059870",
   745 => x"c248c087",
   746 => x"2648c187",
   747 => x"1e4f264b",
   748 => x"4b711e73",
   749 => x"bff0f4c2",
   750 => x"4aa3c449",
   751 => x"8ac24a6a",
   752 => x"bfccf0c2",
   753 => x"49a17292",
   754 => x"bfd0f0c2",
   755 => x"729a6b4a",
   756 => x"fec049a1",
   757 => x"66c859d4",
   758 => x"c4e5711e",
   759 => x"7086c487",
   760 => x"87c40598",
   761 => x"87c248c0",
   762 => x"4b2648c1",
   763 => x"5e0e4f26",
   764 => x"0e5d5c5b",
   765 => x"4b7186e4",
   766 => x"4866ecc0",
   767 => x"a6cc28c9",
   768 => x"d0f0c258",
   769 => x"b9ff49bf",
   770 => x"66c84871",
   771 => x"58a6d498",
   772 => x"986b4871",
   773 => x"c458a6d0",
   774 => x"a6c47ea3",
   775 => x"78bf6e48",
   776 => x"cc4866d0",
   777 => x"c605a866",
   778 => x"7b66c887",
   779 => x"d487c6c3",
   780 => x"ffc148a6",
   781 => x"ffffffff",
   782 => x"ff80c478",
   783 => x"d44ac078",
   784 => x"49724da3",
   785 => x"a17591c8",
   786 => x"4c66d049",
   787 => x"b7c08c69",
   788 => x"87cd04ac",
   789 => x"acb766d4",
   790 => x"dc87c603",
   791 => x"a6d85aa6",
   792 => x"c682c15c",
   793 => x"ff04aab7",
   794 => x"66d887d5",
   795 => x"a8b7c048",
   796 => x"d887d004",
   797 => x"91c84966",
   798 => x"2149a175",
   799 => x"69486e7b",
   800 => x"c087c978",
   801 => x"49a3cc7b",
   802 => x"7869486e",
   803 => x"6b4866c8",
   804 => x"58a6cc88",
   805 => x"bfccf0c2",
   806 => x"7090c848",
   807 => x"4866c87e",
   808 => x"c901a86e",
   809 => x"4866c887",
   810 => x"c003a86e",
   811 => x"c4c187fd",
   812 => x"bf6e7ea3",
   813 => x"7591c849",
   814 => x"66cc49a1",
   815 => x"49bf6e79",
   816 => x"a17591c8",
   817 => x"6681c449",
   818 => x"48a6d079",
   819 => x"d078bf6e",
   820 => x"a8c54866",
   821 => x"c487c705",
   822 => x"78c048a6",
   823 => x"66d087c8",
   824 => x"c880c148",
   825 => x"486e58a6",
   826 => x"c87866c4",
   827 => x"49731e66",
   828 => x"c487f0f8",
   829 => x"cce8c286",
   830 => x"f949731e",
   831 => x"a3d087f2",
   832 => x"66f0c049",
   833 => x"268ee079",
   834 => x"264c264d",
   835 => x"0e4f264b",
   836 => x"0e5c5b5e",
   837 => x"4bc04a71",
   838 => x"c0029a72",
   839 => x"a2da87e0",
   840 => x"4b699f49",
   841 => x"bfd4f0c2",
   842 => x"d487cf02",
   843 => x"699f49a2",
   844 => x"ffc04c49",
   845 => x"34d09cff",
   846 => x"4cc087c2",
   847 => x"9b73b374",
   848 => x"4a87df02",
   849 => x"f0c28ac2",
   850 => x"9249bfcc",
   851 => x"bff0f4c2",
   852 => x"c2807248",
   853 => x"7158d0f5",
   854 => x"c230c448",
   855 => x"c058dcf0",
   856 => x"f4c287e9",
   857 => x"c24bbff4",
   858 => x"c248ccf5",
   859 => x"78bff8f4",
   860 => x"bfd4f0c2",
   861 => x"c287c902",
   862 => x"49bfccf0",
   863 => x"87c731c4",
   864 => x"bffcf4c2",
   865 => x"c231c449",
   866 => x"c259dcf0",
   867 => x"265bccf5",
   868 => x"264b264c",
   869 => x"5b5e0e4f",
   870 => x"f00e5d5c",
   871 => x"59a6c886",
   872 => x"ffffffcf",
   873 => x"7ec04cf8",
   874 => x"d80266c4",
   875 => x"c8e8c287",
   876 => x"c278c048",
   877 => x"c248c0e8",
   878 => x"78bfccf5",
   879 => x"48c4e8c2",
   880 => x"bfc8f5c2",
   881 => x"e9f0c278",
   882 => x"c250c048",
   883 => x"49bfd8f0",
   884 => x"bfc8e8c2",
   885 => x"03aa714a",
   886 => x"7287ccc4",
   887 => x"0599cf49",
   888 => x"c087eac0",
   889 => x"c248d0fe",
   890 => x"78bfc0e8",
   891 => x"1ecce8c2",
   892 => x"bfc0e8c2",
   893 => x"c0e8c249",
   894 => x"78a1c148",
   895 => x"f5dfff71",
   896 => x"c086c487",
   897 => x"c248ccfe",
   898 => x"cc78cce8",
   899 => x"ccfec087",
   900 => x"e0c048bf",
   901 => x"d0fec080",
   902 => x"c8e8c258",
   903 => x"80c148bf",
   904 => x"58cce8c2",
   905 => x"000f8c27",
   906 => x"bf97bf00",
   907 => x"c2029d4d",
   908 => x"e5c387e5",
   909 => x"dec202ad",
   910 => x"ccfec087",
   911 => x"a3cb4bbf",
   912 => x"cf4c1149",
   913 => x"d2c105ac",
   914 => x"df497587",
   915 => x"cd89c199",
   916 => x"dcf0c291",
   917 => x"4aa3c181",
   918 => x"a3c35112",
   919 => x"c551124a",
   920 => x"51124aa3",
   921 => x"124aa3c7",
   922 => x"4aa3c951",
   923 => x"a3ce5112",
   924 => x"d051124a",
   925 => x"51124aa3",
   926 => x"124aa3d2",
   927 => x"4aa3d451",
   928 => x"a3d65112",
   929 => x"d851124a",
   930 => x"51124aa3",
   931 => x"124aa3dc",
   932 => x"4aa3de51",
   933 => x"7ec15112",
   934 => x"7487fcc0",
   935 => x"0599c849",
   936 => x"7487edc0",
   937 => x"0599d049",
   938 => x"e0c087d3",
   939 => x"ccc00266",
   940 => x"c0497387",
   941 => x"700f66e0",
   942 => x"d3c00298",
   943 => x"c0056e87",
   944 => x"f0c287c6",
   945 => x"50c048dc",
   946 => x"bfccfec0",
   947 => x"87e9c248",
   948 => x"48e9f0c2",
   949 => x"c27e50c0",
   950 => x"49bfd8f0",
   951 => x"bfc8e8c2",
   952 => x"04aa714a",
   953 => x"cf87f4fb",
   954 => x"f8ffffff",
   955 => x"ccf5c24c",
   956 => x"c8c005bf",
   957 => x"d4f0c287",
   958 => x"fac102bf",
   959 => x"c4e8c287",
   960 => x"c0eb49bf",
   961 => x"c8e8c287",
   962 => x"48a6c458",
   963 => x"bfc4e8c2",
   964 => x"d4f0c278",
   965 => x"dbc002bf",
   966 => x"4966c487",
   967 => x"a9749974",
   968 => x"87c8c002",
   969 => x"c048a6c8",
   970 => x"87e7c078",
   971 => x"c148a6c8",
   972 => x"87dfc078",
   973 => x"cf4966c4",
   974 => x"a999f8ff",
   975 => x"87c8c002",
   976 => x"c048a6cc",
   977 => x"87c5c078",
   978 => x"c148a6cc",
   979 => x"48a6c878",
   980 => x"c87866cc",
   981 => x"dec00566",
   982 => x"4966c487",
   983 => x"f0c289c2",
   984 => x"c291bfcc",
   985 => x"48bff0f4",
   986 => x"e8c28071",
   987 => x"e8c258c4",
   988 => x"78c048c8",
   989 => x"c087d4f9",
   990 => x"ffffcf48",
   991 => x"f04cf8ff",
   992 => x"264d268e",
   993 => x"264b264c",
   994 => x"0000004f",
   995 => x"00000000",
   996 => x"ffffffff",
   997 => x"48d4ff1e",
   998 => x"6878ffc3",
   999 => x"1e4f2648",
  1000 => x"c348d4ff",
  1001 => x"d0ff78ff",
  1002 => x"78e1c048",
  1003 => x"d448d4ff",
  1004 => x"1e4f2678",
  1005 => x"c048d0ff",
  1006 => x"4f2678e0",
  1007 => x"87d4ff1e",
  1008 => x"02994970",
  1009 => x"fbc087c6",
  1010 => x"87f105a9",
  1011 => x"4f264871",
  1012 => x"5c5b5e0e",
  1013 => x"c04b710e",
  1014 => x"87f8fe4c",
  1015 => x"02994970",
  1016 => x"c087f9c0",
  1017 => x"c002a9ec",
  1018 => x"fbc087f2",
  1019 => x"ebc002a9",
  1020 => x"b766cc87",
  1021 => x"87c703ac",
  1022 => x"c20266d0",
  1023 => x"71537187",
  1024 => x"87c20299",
  1025 => x"cbfe84c1",
  1026 => x"99497087",
  1027 => x"c087cd02",
  1028 => x"c702a9ec",
  1029 => x"a9fbc087",
  1030 => x"87d5ff05",
  1031 => x"c30266d0",
  1032 => x"7b97c087",
  1033 => x"05a9fbc0",
  1034 => x"4a7487c7",
  1035 => x"c28a0ac0",
  1036 => x"724a7487",
  1037 => x"264c2648",
  1038 => x"1e4f264b",
  1039 => x"7087d5fd",
  1040 => x"a9f0c049",
  1041 => x"c087c904",
  1042 => x"c301a9f9",
  1043 => x"89f0c087",
  1044 => x"04a9c1c1",
  1045 => x"dac187c9",
  1046 => x"87c301a9",
  1047 => x"7189f7c0",
  1048 => x"0e4f2648",
  1049 => x"5d5c5b5e",
  1050 => x"7186f80e",
  1051 => x"fc7ec04c",
  1052 => x"4bc087ed",
  1053 => x"97c4c4c1",
  1054 => x"a9c049bf",
  1055 => x"fc87cf04",
  1056 => x"83c187fa",
  1057 => x"97c4c4c1",
  1058 => x"06ab49bf",
  1059 => x"c4c187f1",
  1060 => x"02bf97c4",
  1061 => x"fbfb87cf",
  1062 => x"99497087",
  1063 => x"c087c602",
  1064 => x"f105a9ec",
  1065 => x"fb4bc087",
  1066 => x"4d7087ea",
  1067 => x"c887e5fb",
  1068 => x"dffb58a6",
  1069 => x"c14a7087",
  1070 => x"49a4c883",
  1071 => x"ad496997",
  1072 => x"c987da05",
  1073 => x"699749a4",
  1074 => x"a966c449",
  1075 => x"ca87ce05",
  1076 => x"699749a4",
  1077 => x"c405aa49",
  1078 => x"d07ec187",
  1079 => x"adecc087",
  1080 => x"c087c602",
  1081 => x"c405adfb",
  1082 => x"c14bc087",
  1083 => x"fe026e7e",
  1084 => x"fefa87f5",
  1085 => x"f8487387",
  1086 => x"264d268e",
  1087 => x"264b264c",
  1088 => x"0000004f",
  1089 => x"1e731e00",
  1090 => x"c84bd4ff",
  1091 => x"d0ff4a66",
  1092 => x"78c5c848",
  1093 => x"c148d4ff",
  1094 => x"7b1178d4",
  1095 => x"f9058ac1",
  1096 => x"48d0ff87",
  1097 => x"4b2678c4",
  1098 => x"5e0e4f26",
  1099 => x"0e5d5c5b",
  1100 => x"7e7186f8",
  1101 => x"f5c21e6e",
  1102 => x"ffe349e0",
  1103 => x"7086c487",
  1104 => x"edc40298",
  1105 => x"f4f1c187",
  1106 => x"496e4cbf",
  1107 => x"c887d4fc",
  1108 => x"cac158a6",
  1109 => x"fcfe1ec0",
  1110 => x"86c487f2",
  1111 => x"87c50566",
  1112 => x"c148a6c4",
  1113 => x"48d0ff78",
  1114 => x"d4ff78c5",
  1115 => x"78d5c148",
  1116 => x"c14966c4",
  1117 => x"c131c689",
  1118 => x"bf97ecf1",
  1119 => x"b071484a",
  1120 => x"7808d4ff",
  1121 => x"c448d0ff",
  1122 => x"dcf5c278",
  1123 => x"d049bf97",
  1124 => x"87dd0299",
  1125 => x"d4ff78c5",
  1126 => x"78d6c148",
  1127 => x"d4ff4ac0",
  1128 => x"78ffc348",
  1129 => x"e0c082c1",
  1130 => x"87f204aa",
  1131 => x"c448d0ff",
  1132 => x"48d4ff78",
  1133 => x"ff78ffc3",
  1134 => x"78c548d0",
  1135 => x"c148d4ff",
  1136 => x"78c178d3",
  1137 => x"c448d0ff",
  1138 => x"acb7c078",
  1139 => x"87cbc206",
  1140 => x"bfe8f5c2",
  1141 => x"7e748c4b",
  1142 => x"c1029b73",
  1143 => x"c0c887dd",
  1144 => x"b7c08b4d",
  1145 => x"87c603ab",
  1146 => x"4da3c0c8",
  1147 => x"f5c24bc0",
  1148 => x"49bf97dc",
  1149 => x"cf0299d0",
  1150 => x"c21ec087",
  1151 => x"e549e0f5",
  1152 => x"86c487ee",
  1153 => x"87d84c70",
  1154 => x"1ecce8c2",
  1155 => x"49e0f5c2",
  1156 => x"7087dde5",
  1157 => x"c21e754c",
  1158 => x"fb49cce8",
  1159 => x"86c887e7",
  1160 => x"c5059c74",
  1161 => x"c148c087",
  1162 => x"1ec187ca",
  1163 => x"49e0f5c2",
  1164 => x"c487f0e3",
  1165 => x"059b7386",
  1166 => x"6e87e3fe",
  1167 => x"acb7c04c",
  1168 => x"c287d106",
  1169 => x"c048e0f5",
  1170 => x"c080d078",
  1171 => x"c280f478",
  1172 => x"78bfecf5",
  1173 => x"01acb7c0",
  1174 => x"ff87f5fd",
  1175 => x"78c548d0",
  1176 => x"c148d4ff",
  1177 => x"78c078d3",
  1178 => x"c448d0ff",
  1179 => x"c048c178",
  1180 => x"48c087c2",
  1181 => x"4d268ef8",
  1182 => x"4b264c26",
  1183 => x"00004f26",
  1184 => x"20746f47",
  1185 => x"69747865",
  1186 => x"0000646e",
  1187 => x"64616f4c",
  1188 => x"2e676e69",
  1189 => x"00002e2e",
  1190 => x"61422080",
  1191 => x"00006b63",
  1192 => x"64616f4c",
  1193 => x"202e2a20",
  1194 => x"00000000",
  1195 => x"0000203a",
  1196 => x"61422080",
  1197 => x"00006b63",
  1198 => x"78452080",
  1199 => x"00007469",
  1200 => x"49204453",
  1201 => x"2e74696e",
  1202 => x"0000002e",
  1203 => x"00004b4f",
  1204 => x"544f4f42",
  1205 => x"20202020",
  1206 => x"004d4f52",
  1207 => x"5c5b5e0e",
  1208 => x"86fc0e5d",
  1209 => x"4bc04d71",
  1210 => x"c004ad4c",
  1211 => x"c1c187e8",
  1212 => x"9c741ee3",
  1213 => x"c087c402",
  1214 => x"c187c24a",
  1215 => x"ea49724a",
  1216 => x"86c487d3",
  1217 => x"83c17e70",
  1218 => x"87c2056e",
  1219 => x"84c14b75",
  1220 => x"ff06ab75",
  1221 => x"486e87d8",
  1222 => x"4d268efc",
  1223 => x"4b264c26",
  1224 => x"5e0e4f26",
  1225 => x"710e5c5b",
  1226 => x"0266cc4b",
  1227 => x"c04c87d8",
  1228 => x"d8028cf0",
  1229 => x"c14a7487",
  1230 => x"87d1028a",
  1231 => x"87cd028a",
  1232 => x"87c9028a",
  1233 => x"497387d9",
  1234 => x"d287dff7",
  1235 => x"c01e7487",
  1236 => x"dbd7c149",
  1237 => x"731e7487",
  1238 => x"d3d7c149",
  1239 => x"2686c887",
  1240 => x"264b264c",
  1241 => x"5b5e0e4f",
  1242 => x"fc0e5d5c",
  1243 => x"494c7186",
  1244 => x"f7c291de",
  1245 => x"85714dc0",
  1246 => x"c1026d97",
  1247 => x"f6c287db",
  1248 => x"7449bff0",
  1249 => x"d3fd7181",
  1250 => x"487e7087",
  1251 => x"f2c00298",
  1252 => x"f4f6c287",
  1253 => x"cb4a704b",
  1254 => x"c5fafe49",
  1255 => x"cc4b7487",
  1256 => x"f8f1c193",
  1257 => x"c183c483",
  1258 => x"747bccca",
  1259 => x"cbc1c149",
  1260 => x"c17b7587",
  1261 => x"bf97f0f1",
  1262 => x"f6c21e49",
  1263 => x"e1fd49f4",
  1264 => x"7486c487",
  1265 => x"f3c0c149",
  1266 => x"c149c087",
  1267 => x"c287cec2",
  1268 => x"c048d8f5",
  1269 => x"e4df4950",
  1270 => x"268efc87",
  1271 => x"264c264d",
  1272 => x"1e4f264b",
  1273 => x"4b711e73",
  1274 => x"f0f6c249",
  1275 => x"fb7181bf",
  1276 => x"4a7087ea",
  1277 => x"87c4029a",
  1278 => x"87d3e449",
  1279 => x"48f0f6c2",
  1280 => x"497378c0",
  1281 => x"2687fac1",
  1282 => x"1e4f264b",
  1283 => x"4b711e73",
  1284 => x"024aa3c4",
  1285 => x"c187d0c1",
  1286 => x"87dc028a",
  1287 => x"f2c0028a",
  1288 => x"c1058a87",
  1289 => x"f6c287d3",
  1290 => x"c102bff0",
  1291 => x"c14887cb",
  1292 => x"f4f6c288",
  1293 => x"87c1c158",
  1294 => x"bff0f6c2",
  1295 => x"c289c649",
  1296 => x"c059f4f6",
  1297 => x"c003a9b7",
  1298 => x"f6c287ef",
  1299 => x"78c048f0",
  1300 => x"c287e6c0",
  1301 => x"02bfecf6",
  1302 => x"f6c287df",
  1303 => x"c148bff0",
  1304 => x"f4f6c280",
  1305 => x"c287d258",
  1306 => x"02bfecf6",
  1307 => x"f6c287cb",
  1308 => x"c648bff0",
  1309 => x"f4f6c280",
  1310 => x"c4497358",
  1311 => x"264b2687",
  1312 => x"5b5e0e4f",
  1313 => x"f00e5d5c",
  1314 => x"59a6d086",
  1315 => x"4dcce8c2",
  1316 => x"f6c24cc0",
  1317 => x"78c148ec",
  1318 => x"c048a6c8",
  1319 => x"c27e7578",
  1320 => x"48bff0f6",
  1321 => x"c106a8c0",
  1322 => x"a6c887c0",
  1323 => x"c27e755c",
  1324 => x"9848cce8",
  1325 => x"87f2c002",
  1326 => x"c14d66c4",
  1327 => x"cc1ee3c1",
  1328 => x"87c40266",
  1329 => x"87c24cc0",
  1330 => x"49744cc1",
  1331 => x"c487c6e3",
  1332 => x"c17e7086",
  1333 => x"4866c885",
  1334 => x"a6cc80c1",
  1335 => x"f0f6c258",
  1336 => x"c503adbf",
  1337 => x"ff056e87",
  1338 => x"4d6e87d1",
  1339 => x"9d754cc0",
  1340 => x"87dcc302",
  1341 => x"1ee3c1c1",
  1342 => x"c70266cc",
  1343 => x"48a6c887",
  1344 => x"87c578c0",
  1345 => x"c148a6c8",
  1346 => x"4966c878",
  1347 => x"c487c6e2",
  1348 => x"487e7086",
  1349 => x"e4c20298",
  1350 => x"81cb4987",
  1351 => x"d0496997",
  1352 => x"d4c10299",
  1353 => x"cc497487",
  1354 => x"f8f1c191",
  1355 => x"e3cfc181",
  1356 => x"c381c879",
  1357 => x"497451ff",
  1358 => x"f7c291de",
  1359 => x"85714dc0",
  1360 => x"7d97c1c2",
  1361 => x"c049a5c1",
  1362 => x"f0c251e0",
  1363 => x"02bf97dc",
  1364 => x"84c187d2",
  1365 => x"c24ba5c2",
  1366 => x"db4adcf0",
  1367 => x"c1f3fe49",
  1368 => x"87d9c187",
  1369 => x"c049a5cd",
  1370 => x"c284c151",
  1371 => x"4a6e4ba5",
  1372 => x"f2fe49cb",
  1373 => x"c4c187ec",
  1374 => x"cc497487",
  1375 => x"f8f1c191",
  1376 => x"e5cdc181",
  1377 => x"dcf0c279",
  1378 => x"d802bf97",
  1379 => x"de497487",
  1380 => x"c284c191",
  1381 => x"714bc0f7",
  1382 => x"dcf0c283",
  1383 => x"fe49dd4a",
  1384 => x"d887fff1",
  1385 => x"de4b7487",
  1386 => x"c0f7c293",
  1387 => x"49a3cb83",
  1388 => x"84c151c0",
  1389 => x"cb4a6e73",
  1390 => x"e5f1fe49",
  1391 => x"4866c887",
  1392 => x"a6cc80c1",
  1393 => x"03acc758",
  1394 => x"6e87c5c0",
  1395 => x"87e4fc05",
  1396 => x"c003acc7",
  1397 => x"f6c287e4",
  1398 => x"78c048ec",
  1399 => x"91cc4974",
  1400 => x"81f8f1c1",
  1401 => x"79e5cdc1",
  1402 => x"91de4974",
  1403 => x"81c0f7c2",
  1404 => x"84c151c0",
  1405 => x"ff04acc7",
  1406 => x"f3c187dc",
  1407 => x"50c048d4",
  1408 => x"d9c180f7",
  1409 => x"cac140d9",
  1410 => x"80c878d8",
  1411 => x"78cbd0c1",
  1412 => x"c04966cc",
  1413 => x"f087e5f7",
  1414 => x"264d268e",
  1415 => x"264b264c",
  1416 => x"1e731e4f",
  1417 => x"cc494b71",
  1418 => x"f8f1c191",
  1419 => x"4aa1c881",
  1420 => x"48ecf1c1",
  1421 => x"a1c95012",
  1422 => x"c4c4c14a",
  1423 => x"ca501248",
  1424 => x"f0f1c181",
  1425 => x"73501148",
  1426 => x"87f5f849",
  1427 => x"4f264b26",
  1428 => x"c049c01e",
  1429 => x"2687c6f8",
  1430 => x"4a711e4f",
  1431 => x"c191cc49",
  1432 => x"c881f8f1",
  1433 => x"d8f5c281",
  1434 => x"c0501148",
  1435 => x"fe49a2f0",
  1436 => x"c087fbec",
  1437 => x"87c5d549",
  1438 => x"ff1e4f26",
  1439 => x"ffc34ad4",
  1440 => x"48d0ff7a",
  1441 => x"de78e1c0",
  1442 => x"487a717a",
  1443 => x"7028b7c8",
  1444 => x"d048717a",
  1445 => x"7a7028b7",
  1446 => x"b7d84871",
  1447 => x"ff7a7028",
  1448 => x"e0c048d0",
  1449 => x"0e4f2678",
  1450 => x"5d5c5b5e",
  1451 => x"7186f40e",
  1452 => x"91cc494d",
  1453 => x"81f8f1c1",
  1454 => x"ca4aa1c8",
  1455 => x"a6c47ea1",
  1456 => x"d4f5c248",
  1457 => x"976e78bf",
  1458 => x"66c44bbf",
  1459 => x"122c734c",
  1460 => x"58a6cc48",
  1461 => x"84c19c70",
  1462 => x"699781c9",
  1463 => x"04acb749",
  1464 => x"4cc087c2",
  1465 => x"4abf976e",
  1466 => x"724966c8",
  1467 => x"c4b9ff31",
  1468 => x"48749966",
  1469 => x"4a703072",
  1470 => x"d8f5c2b1",
  1471 => x"f9fd7159",
  1472 => x"c21ec787",
  1473 => x"1ebfe8f6",
  1474 => x"1ef8f1c1",
  1475 => x"97d8f5c2",
  1476 => x"f4c149bf",
  1477 => x"c0497587",
  1478 => x"e887e1f3",
  1479 => x"264d268e",
  1480 => x"264b264c",
  1481 => x"1e731e4f",
  1482 => x"fd494b71",
  1483 => x"497387f9",
  1484 => x"2687f4fd",
  1485 => x"1e4f264b",
  1486 => x"4b711e73",
  1487 => x"024aa3c2",
  1488 => x"8ac187d6",
  1489 => x"87e2c005",
  1490 => x"bfe8f6c2",
  1491 => x"4887db02",
  1492 => x"f6c288c1",
  1493 => x"87d258ec",
  1494 => x"bfecf6c2",
  1495 => x"c287cb02",
  1496 => x"48bfe8f6",
  1497 => x"f6c280c1",
  1498 => x"1ec758ec",
  1499 => x"bfe8f6c2",
  1500 => x"f8f1c11e",
  1501 => x"d8f5c21e",
  1502 => x"cc49bf97",
  1503 => x"c0497387",
  1504 => x"f487f9f1",
  1505 => x"264b268e",
  1506 => x"5b5e0e4f",
  1507 => x"ff0e5d5c",
  1508 => x"e8c086cc",
  1509 => x"a6cc59a6",
  1510 => x"c478c048",
  1511 => x"c478c080",
  1512 => x"c478c080",
  1513 => x"66c8c180",
  1514 => x"c180c478",
  1515 => x"c180c478",
  1516 => x"ecf6c278",
  1517 => x"ff78c148",
  1518 => x"ff87e4df",
  1519 => x"ff87fddf",
  1520 => x"7087d1df",
  1521 => x"adfbc04d",
  1522 => x"87f3c102",
  1523 => x"0566e4c0",
  1524 => x"c187e8c1",
  1525 => x"c44a66c4",
  1526 => x"c17e6a82",
  1527 => x"6e48e0ca",
  1528 => x"20412049",
  1529 => x"c1511041",
  1530 => x"c14866c4",
  1531 => x"6a78e1d8",
  1532 => x"7581c749",
  1533 => x"66c4c151",
  1534 => x"c181c849",
  1535 => x"48a6dc51",
  1536 => x"c4c178c2",
  1537 => x"81c94966",
  1538 => x"c4c151c0",
  1539 => x"81ca4966",
  1540 => x"1ec151c0",
  1541 => x"496a1ed8",
  1542 => x"deff81c8",
  1543 => x"86c887f2",
  1544 => x"4866c8c1",
  1545 => x"c701a8c0",
  1546 => x"48a6d487",
  1547 => x"87cf78c1",
  1548 => x"4866c8c1",
  1549 => x"a6dc88c1",
  1550 => x"ff87c458",
  1551 => x"7587fddd",
  1552 => x"f2cb029d",
  1553 => x"4866d487",
  1554 => x"a866ccc1",
  1555 => x"87e7cb03",
  1556 => x"dcff7ec0",
  1557 => x"4d7087fe",
  1558 => x"88c6c148",
  1559 => x"7058a6c8",
  1560 => x"d6c10298",
  1561 => x"88c94887",
  1562 => x"7058a6c8",
  1563 => x"d8c50298",
  1564 => x"88c14887",
  1565 => x"7058a6c8",
  1566 => x"f8c20298",
  1567 => x"88c34887",
  1568 => x"7058a6c8",
  1569 => x"87cf0298",
  1570 => x"c888c148",
  1571 => x"987058a6",
  1572 => x"87f5c402",
  1573 => x"c087ffc9",
  1574 => x"dbff7ef0",
  1575 => x"4d7087f6",
  1576 => x"02adecc0",
  1577 => x"7e7587c2",
  1578 => x"02adecc0",
  1579 => x"dbff87cd",
  1580 => x"4d7087e2",
  1581 => x"05adecc0",
  1582 => x"c087f3ff",
  1583 => x"c10566e4",
  1584 => x"ecc087ea",
  1585 => x"87c402ad",
  1586 => x"87c8dbff",
  1587 => x"1eca1ec0",
  1588 => x"cc4b66dc",
  1589 => x"66ccc193",
  1590 => x"4ca3c483",
  1591 => x"dbff496c",
  1592 => x"1ec187ee",
  1593 => x"496c1ede",
  1594 => x"87e4dbff",
  1595 => x"d8c186d0",
  1596 => x"a3c87be1",
  1597 => x"5166dc49",
  1598 => x"c049a3c9",
  1599 => x"ca5166e0",
  1600 => x"516e49a3",
  1601 => x"c14866dc",
  1602 => x"a6e0c080",
  1603 => x"4866d458",
  1604 => x"04a866d8",
  1605 => x"66d487cb",
  1606 => x"d880c148",
  1607 => x"fbc758a6",
  1608 => x"4866d887",
  1609 => x"a6dc88c1",
  1610 => x"87f0c758",
  1611 => x"87ccdaff",
  1612 => x"e7c74d70",
  1613 => x"c2dcff87",
  1614 => x"58a6d087",
  1615 => x"06a866d0",
  1616 => x"d087c6c0",
  1617 => x"66cc48a6",
  1618 => x"eedbff78",
  1619 => x"a8ecc087",
  1620 => x"87f5c105",
  1621 => x"0566e4c0",
  1622 => x"d487e5c1",
  1623 => x"91cc4966",
  1624 => x"8166c4c1",
  1625 => x"6a4aa1c4",
  1626 => x"4aa1c84c",
  1627 => x"c15266cc",
  1628 => x"ff79d9d9",
  1629 => x"7087ddd8",
  1630 => x"da029d4d",
  1631 => x"adfbc087",
  1632 => x"7587d402",
  1633 => x"cbd8ff54",
  1634 => x"9d4d7087",
  1635 => x"87c7c002",
  1636 => x"05adfbc0",
  1637 => x"c087ecff",
  1638 => x"c1c254e0",
  1639 => x"7c97c054",
  1640 => x"d84866d4",
  1641 => x"c004a866",
  1642 => x"66d487cb",
  1643 => x"d880c148",
  1644 => x"e7c558a6",
  1645 => x"4866d887",
  1646 => x"a6dc88c1",
  1647 => x"87dcc558",
  1648 => x"87f8d7ff",
  1649 => x"d3c54d70",
  1650 => x"4866cc87",
  1651 => x"a866e4c0",
  1652 => x"87f4c405",
  1653 => x"48a6e8c0",
  1654 => x"d9ff78c0",
  1655 => x"7e7087dd",
  1656 => x"87d7d9ff",
  1657 => x"58a6f0c0",
  1658 => x"05a8ecc0",
  1659 => x"a687c7c0",
  1660 => x"c0786e48",
  1661 => x"d6ff87c4",
  1662 => x"66d487da",
  1663 => x"c191cc49",
  1664 => x"714866c4",
  1665 => x"58a6c880",
  1666 => x"c84a66c4",
  1667 => x"4966c482",
  1668 => x"516e81ca",
  1669 => x"4966ecc0",
  1670 => x"896e81c1",
  1671 => x"307148c1",
  1672 => x"89c14970",
  1673 => x"c27a9771",
  1674 => x"49bfd4f5",
  1675 => x"6a97296e",
  1676 => x"9871484a",
  1677 => x"58a6f4c0",
  1678 => x"c44866c4",
  1679 => x"58a6cc80",
  1680 => x"4cbf66c8",
  1681 => x"4866e4c0",
  1682 => x"02a866cc",
  1683 => x"c087c5c0",
  1684 => x"87c2c07e",
  1685 => x"1e6e7ec1",
  1686 => x"741ee0c0",
  1687 => x"efd5ff49",
  1688 => x"7086c887",
  1689 => x"adb7c04d",
  1690 => x"87d4c106",
  1691 => x"66c88475",
  1692 => x"e0c049bf",
  1693 => x"4b897481",
  1694 => x"4aeccac1",
  1695 => x"e1defe71",
  1696 => x"7484c287",
  1697 => x"66e8c07e",
  1698 => x"c080c148",
  1699 => x"c058a6ec",
  1700 => x"c14966f0",
  1701 => x"02a97081",
  1702 => x"c087c5c0",
  1703 => x"87c2c04c",
  1704 => x"1e744cc1",
  1705 => x"49bf66cc",
  1706 => x"c481e0c0",
  1707 => x"1e718966",
  1708 => x"ff4966c8",
  1709 => x"c887d9d4",
  1710 => x"a8b7c086",
  1711 => x"87c5ff01",
  1712 => x"0266e8c0",
  1713 => x"c487d3c0",
  1714 => x"81c94966",
  1715 => x"5166e8c0",
  1716 => x"c14866c4",
  1717 => x"c078e7da",
  1718 => x"66c487ce",
  1719 => x"c281c949",
  1720 => x"4866c451",
  1721 => x"78e5dcc1",
  1722 => x"d84866d4",
  1723 => x"c004a866",
  1724 => x"66d487cb",
  1725 => x"d880c148",
  1726 => x"d1c058a6",
  1727 => x"4866d887",
  1728 => x"a6dc88c1",
  1729 => x"87c6c058",
  1730 => x"87f0d2ff",
  1731 => x"a6cc4d70",
  1732 => x"c078c048",
  1733 => x"d2ff87c6",
  1734 => x"4d7087e2",
  1735 => x"4866e0c0",
  1736 => x"e4c080c1",
  1737 => x"9d7558a6",
  1738 => x"87cbc002",
  1739 => x"c14866d4",
  1740 => x"04a866cc",
  1741 => x"d487d9f4",
  1742 => x"a8c74866",
  1743 => x"87e1c003",
  1744 => x"c24c66d4",
  1745 => x"c048ecf6",
  1746 => x"cc497478",
  1747 => x"66c4c191",
  1748 => x"4aa1c481",
  1749 => x"52c04a6a",
  1750 => x"c784c179",
  1751 => x"e2ff04ac",
  1752 => x"66e4c087",
  1753 => x"87e2c002",
  1754 => x"4966c4c1",
  1755 => x"c181d4c1",
  1756 => x"c14a66c4",
  1757 => x"52c082dc",
  1758 => x"79d9d9c1",
  1759 => x"4966c4c1",
  1760 => x"c181d8c1",
  1761 => x"c079f0ca",
  1762 => x"c4c187d6",
  1763 => x"d4c14966",
  1764 => x"66c4c181",
  1765 => x"82d8c14a",
  1766 => x"7af8cac1",
  1767 => x"79d0d9c1",
  1768 => x"4966c4c1",
  1769 => x"c181e0c1",
  1770 => x"ff79f7dc",
  1771 => x"d087c4d0",
  1772 => x"ccff4866",
  1773 => x"264d268e",
  1774 => x"264b264c",
  1775 => x"1ec71e4f",
  1776 => x"bfe8f6c2",
  1777 => x"f8f1c11e",
  1778 => x"d8f5c21e",
  1779 => x"ee49bf97",
  1780 => x"f1c187f7",
  1781 => x"e1c049f8",
  1782 => x"8ef487f0",
  1783 => x"c11e4f26",
  1784 => x"c048ecf1",
  1785 => x"e4f3c150",
  1786 => x"d4ff49bf",
  1787 => x"48c087fc",
  1788 => x"731e4f26",
  1789 => x"87cec71e",
  1790 => x"48f4f6c2",
  1791 => x"d4ff50c0",
  1792 => x"78ffc348",
  1793 => x"49c0cbc1",
  1794 => x"87fdd6fe",
  1795 => x"87d0e2fe",
  1796 => x"cd029870",
  1797 => x"eeebfe87",
  1798 => x"02987087",
  1799 => x"4ac187c4",
  1800 => x"4ac087c2",
  1801 => x"c8029a72",
  1802 => x"cccbc187",
  1803 => x"d8d6fe49",
  1804 => x"e8f6c287",
  1805 => x"c278c048",
  1806 => x"c048d8f5",
  1807 => x"fcfd4950",
  1808 => x"87dafe87",
  1809 => x"029b4b70",
  1810 => x"f3c187cf",
  1811 => x"49c75bd4",
  1812 => x"c187e9de",
  1813 => x"c4e0c049",
  1814 => x"87f3c287",
  1815 => x"87cae1c0",
  1816 => x"87dcefc0",
  1817 => x"2687f5ff",
  1818 => x"004f264b",
  1819 => x"00000000",
  1820 => x"00000000",
  1821 => x"00000001",
  1822 => x"00001365",
  1823 => x"00002dc0",
  1824 => x"94000000",
  1825 => x"00001365",
  1826 => x"00002dde",
  1827 => x"94000000",
  1828 => x"00001365",
  1829 => x"00002dfc",
  1830 => x"94000000",
  1831 => x"00001365",
  1832 => x"00002e1a",
  1833 => x"94000000",
  1834 => x"00001365",
  1835 => x"00002e38",
  1836 => x"94000000",
  1837 => x"00001365",
  1838 => x"00002e56",
  1839 => x"94000000",
  1840 => x"00001365",
  1841 => x"00002e74",
  1842 => x"94000000",
  1843 => x"00001659",
  1844 => x"00000000",
  1845 => x"94000000",
  1846 => x"0000140b",
  1847 => x"00000000",
  1848 => x"94000000",
  1849 => x"000012d0",
  1850 => x"db86fc1e",
  1851 => x"fc7e7087",
  1852 => x"1e4f268e",
  1853 => x"c048f0fe",
  1854 => x"7909cd78",
  1855 => x"1e4f2609",
  1856 => x"49e8f3c1",
  1857 => x"4f2687ed",
  1858 => x"bff0fe1e",
  1859 => x"1e4f2648",
  1860 => x"c148f0fe",
  1861 => x"1e4f2678",
  1862 => x"c048f0fe",
  1863 => x"1e4f2678",
  1864 => x"52c04a71",
  1865 => x"0e4f2651",
  1866 => x"5d5c5b5e",
  1867 => x"7186f40e",
  1868 => x"7e6d974d",
  1869 => x"974ca5c1",
  1870 => x"a6c8486c",
  1871 => x"c4486e58",
  1872 => x"c505a866",
  1873 => x"c048ff87",
  1874 => x"caff87e6",
  1875 => x"49a5c287",
  1876 => x"714b6c97",
  1877 => x"6b974ba3",
  1878 => x"7e6c974b",
  1879 => x"80c1486e",
  1880 => x"c758a6c8",
  1881 => x"58a6cc98",
  1882 => x"fe7c9770",
  1883 => x"487387e1",
  1884 => x"4d268ef4",
  1885 => x"4b264c26",
  1886 => x"731e4f26",
  1887 => x"fe86f41e",
  1888 => x"bfe087d5",
  1889 => x"e0c0494b",
  1890 => x"c00299c0",
  1891 => x"4a7387ea",
  1892 => x"c29affc3",
  1893 => x"bf97e8fa",
  1894 => x"eafac249",
  1895 => x"c2517281",
  1896 => x"bf97e8fa",
  1897 => x"c1486e7e",
  1898 => x"58a6c880",
  1899 => x"a6cc98c7",
  1900 => x"e8fac258",
  1901 => x"5066c848",
  1902 => x"7087cdfd",
  1903 => x"87cffd7e",
  1904 => x"4b268ef4",
  1905 => x"c21e4f26",
  1906 => x"fd49e8fa",
  1907 => x"f5c187d1",
  1908 => x"defc49fa",
  1909 => x"87e8c487",
  1910 => x"5e0e4f26",
  1911 => x"0e5d5c5b",
  1912 => x"7e7186fc",
  1913 => x"c24dd4ff",
  1914 => x"fc49e8fa",
  1915 => x"4b7087f9",
  1916 => x"04abb7c0",
  1917 => x"c387f5c2",
  1918 => x"c905abf0",
  1919 => x"f8fac187",
  1920 => x"c278c148",
  1921 => x"e0c387d6",
  1922 => x"87c905ab",
  1923 => x"48fcfac1",
  1924 => x"c7c278c1",
  1925 => x"fcfac187",
  1926 => x"87c602bf",
  1927 => x"4ca3c0c2",
  1928 => x"4c7387c2",
  1929 => x"bff8fac1",
  1930 => x"87e0c002",
  1931 => x"b7c44974",
  1932 => x"fbc19129",
  1933 => x"4a7481c0",
  1934 => x"92c29acf",
  1935 => x"307248c1",
  1936 => x"baff4a70",
  1937 => x"98694872",
  1938 => x"87db7970",
  1939 => x"b7c44974",
  1940 => x"fbc19129",
  1941 => x"4a7481c0",
  1942 => x"92c29acf",
  1943 => x"307248c3",
  1944 => x"69484a70",
  1945 => x"6e7970b0",
  1946 => x"87e4c005",
  1947 => x"c848d0ff",
  1948 => x"7dc578e1",
  1949 => x"bffcfac1",
  1950 => x"c387c302",
  1951 => x"fac17de0",
  1952 => x"c302bff8",
  1953 => x"7df0c387",
  1954 => x"d0ff7d73",
  1955 => x"78e0c048",
  1956 => x"48fcfac1",
  1957 => x"fac178c0",
  1958 => x"78c048f8",
  1959 => x"49e8fac2",
  1960 => x"7087c4fa",
  1961 => x"abb7c04b",
  1962 => x"87cbfd03",
  1963 => x"8efc48c0",
  1964 => x"4c264d26",
  1965 => x"4f264b26",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"84848484",
  1970 => x"84848484",
  1971 => x"84848484",
  1972 => x"84848484",
  1973 => x"84848484",
  1974 => x"84848484",
  1975 => x"84848484",
  1976 => x"84848484",
  1977 => x"84848484",
  1978 => x"84848484",
  1979 => x"84848484",
  1980 => x"84848484",
  1981 => x"84848484",
  1982 => x"84848484",
  1983 => x"84848484",
  1984 => x"724ac01e",
  1985 => x"c191c449",
  1986 => x"c081c0fb",
  1987 => x"d082c179",
  1988 => x"ee04aab7",
  1989 => x"0e4f2687",
  1990 => x"5d5c5b5e",
  1991 => x"f74d710e",
  1992 => x"4a7587f5",
  1993 => x"922ab7c4",
  1994 => x"82c0fbc1",
  1995 => x"9ccf4c75",
  1996 => x"496a94c2",
  1997 => x"c32b744b",
  1998 => x"7448c29b",
  1999 => x"ff4c7030",
  2000 => x"714874bc",
  2001 => x"f77a7098",
  2002 => x"487387c5",
  2003 => x"4c264d26",
  2004 => x"4f264b26",
  2005 => x"48d0ff1e",
  2006 => x"7178e1c8",
  2007 => x"08d4ff48",
  2008 => x"1e4f2678",
  2009 => x"c848d0ff",
  2010 => x"487178e1",
  2011 => x"7808d4ff",
  2012 => x"ff4866c4",
  2013 => x"267808d4",
  2014 => x"4a711e4f",
  2015 => x"1e4966c4",
  2016 => x"deff4972",
  2017 => x"48d0ff87",
  2018 => x"fc78e0c0",
  2019 => x"1e4f268e",
  2020 => x"4b711e73",
  2021 => x"1e4966c8",
  2022 => x"e0c14a73",
  2023 => x"d8ff49a2",
  2024 => x"268efc87",
  2025 => x"1e4f264b",
  2026 => x"c848d0ff",
  2027 => x"487178c9",
  2028 => x"7808d4ff",
  2029 => x"711e4f26",
  2030 => x"87eb494a",
  2031 => x"c848d0ff",
  2032 => x"1e4f2678",
  2033 => x"4b711e73",
  2034 => x"bfc0fbc2",
  2035 => x"c287c302",
  2036 => x"d0ff87eb",
  2037 => x"78c9c848",
  2038 => x"e0c04873",
  2039 => x"08d4ffb0",
  2040 => x"f4fac278",
  2041 => x"c878c048",
  2042 => x"87c50266",
  2043 => x"c249ffc3",
  2044 => x"c249c087",
  2045 => x"cc59fcfa",
  2046 => x"87c60266",
  2047 => x"4ad5d5c5",
  2048 => x"ffcf87c4",
  2049 => x"fbc24aff",
  2050 => x"fbc25ac0",
  2051 => x"78c148c0",
  2052 => x"4f264b26",
  2053 => x"5c5b5e0e",
  2054 => x"4d710e5d",
  2055 => x"bffcfac2",
  2056 => x"029d754b",
  2057 => x"c84987cb",
  2058 => x"fcfec191",
  2059 => x"c482714a",
  2060 => x"fcc2c287",
  2061 => x"124cc04a",
  2062 => x"c2997349",
  2063 => x"48bff8fa",
  2064 => x"d4ffb871",
  2065 => x"b7c17808",
  2066 => x"b7c8842b",
  2067 => x"87e704ac",
  2068 => x"bff4fac2",
  2069 => x"c280c848",
  2070 => x"2658f8fa",
  2071 => x"264c264d",
  2072 => x"1e4f264b",
  2073 => x"4b711e73",
  2074 => x"029a4a13",
  2075 => x"497287cb",
  2076 => x"1387e1fe",
  2077 => x"f5059a4a",
  2078 => x"264b2687",
  2079 => x"fac21e4f",
  2080 => x"c249bff4",
  2081 => x"c148f4fa",
  2082 => x"c0c478a1",
  2083 => x"db03a9b7",
  2084 => x"48d4ff87",
  2085 => x"bff8fac2",
  2086 => x"f4fac278",
  2087 => x"fac249bf",
  2088 => x"a1c148f4",
  2089 => x"b7c0c478",
  2090 => x"87e504a9",
  2091 => x"c848d0ff",
  2092 => x"c0fbc278",
  2093 => x"2678c048",
  2094 => x"0000004f",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"5f000000",
  2098 => x"0000005f",
  2099 => x"00030300",
  2100 => x"00000303",
  2101 => x"147f7f14",
  2102 => x"00147f7f",
  2103 => x"6b2e2400",
  2104 => x"00123a6b",
  2105 => x"18366a4c",
  2106 => x"0032566c",
  2107 => x"594f7e30",
  2108 => x"40683a77",
  2109 => x"07040000",
  2110 => x"00000003",
  2111 => x"3e1c0000",
  2112 => x"00004163",
  2113 => x"63410000",
  2114 => x"00001c3e",
  2115 => x"1c3e2a08",
  2116 => x"082a3e1c",
  2117 => x"3e080800",
  2118 => x"0008083e",
  2119 => x"e0800000",
  2120 => x"00000060",
  2121 => x"08080800",
  2122 => x"00080808",
  2123 => x"60000000",
  2124 => x"00000060",
  2125 => x"18306040",
  2126 => x"0103060c",
  2127 => x"597f3e00",
  2128 => x"003e7f4d",
  2129 => x"7f060400",
  2130 => x"0000007f",
  2131 => x"71634200",
  2132 => x"00464f59",
  2133 => x"49632200",
  2134 => x"00367f49",
  2135 => x"13161c18",
  2136 => x"00107f7f",
  2137 => x"45672700",
  2138 => x"00397d45",
  2139 => x"4b7e3c00",
  2140 => x"00307949",
  2141 => x"71010100",
  2142 => x"00070f79",
  2143 => x"497f3600",
  2144 => x"00367f49",
  2145 => x"494f0600",
  2146 => x"001e3f69",
  2147 => x"66000000",
  2148 => x"00000066",
  2149 => x"e6800000",
  2150 => x"00000066",
  2151 => x"14080800",
  2152 => x"00222214",
  2153 => x"14141400",
  2154 => x"00141414",
  2155 => x"14222200",
  2156 => x"00080814",
  2157 => x"51030200",
  2158 => x"00060f59",
  2159 => x"5d417f3e",
  2160 => x"001e1f55",
  2161 => x"097f7e00",
  2162 => x"007e7f09",
  2163 => x"497f7f00",
  2164 => x"00367f49",
  2165 => x"633e1c00",
  2166 => x"00414141",
  2167 => x"417f7f00",
  2168 => x"001c3e63",
  2169 => x"497f7f00",
  2170 => x"00414149",
  2171 => x"097f7f00",
  2172 => x"00010109",
  2173 => x"417f3e00",
  2174 => x"007a7b49",
  2175 => x"087f7f00",
  2176 => x"007f7f08",
  2177 => x"7f410000",
  2178 => x"0000417f",
  2179 => x"40602000",
  2180 => x"003f7f40",
  2181 => x"1c087f7f",
  2182 => x"00416336",
  2183 => x"407f7f00",
  2184 => x"00404040",
  2185 => x"0c067f7f",
  2186 => x"007f7f06",
  2187 => x"0c067f7f",
  2188 => x"007f7f18",
  2189 => x"417f3e00",
  2190 => x"003e7f41",
  2191 => x"097f7f00",
  2192 => x"00060f09",
  2193 => x"61417f3e",
  2194 => x"00407e7f",
  2195 => x"097f7f00",
  2196 => x"00667f19",
  2197 => x"4d6f2600",
  2198 => x"00327b59",
  2199 => x"7f010100",
  2200 => x"0001017f",
  2201 => x"407f3f00",
  2202 => x"003f7f40",
  2203 => x"703f0f00",
  2204 => x"000f3f70",
  2205 => x"18307f7f",
  2206 => x"007f7f30",
  2207 => x"1c366341",
  2208 => x"4163361c",
  2209 => x"7c060301",
  2210 => x"0103067c",
  2211 => x"4d597161",
  2212 => x"00414347",
  2213 => x"7f7f0000",
  2214 => x"00004141",
  2215 => x"0c060301",
  2216 => x"40603018",
  2217 => x"41410000",
  2218 => x"00007f7f",
  2219 => x"03060c08",
  2220 => x"00080c06",
  2221 => x"80808080",
  2222 => x"00808080",
  2223 => x"03000000",
  2224 => x"00000407",
  2225 => x"54742000",
  2226 => x"00787c54",
  2227 => x"447f7f00",
  2228 => x"00387c44",
  2229 => x"447c3800",
  2230 => x"00004444",
  2231 => x"447c3800",
  2232 => x"007f7f44",
  2233 => x"547c3800",
  2234 => x"00185c54",
  2235 => x"7f7e0400",
  2236 => x"00000505",
  2237 => x"a4bc1800",
  2238 => x"007cfca4",
  2239 => x"047f7f00",
  2240 => x"00787c04",
  2241 => x"3d000000",
  2242 => x"0000407d",
  2243 => x"80808000",
  2244 => x"00007dfd",
  2245 => x"107f7f00",
  2246 => x"00446c38",
  2247 => x"3f000000",
  2248 => x"0000407f",
  2249 => x"180c7c7c",
  2250 => x"00787c0c",
  2251 => x"047c7c00",
  2252 => x"00787c04",
  2253 => x"447c3800",
  2254 => x"00387c44",
  2255 => x"24fcfc00",
  2256 => x"00183c24",
  2257 => x"243c1800",
  2258 => x"00fcfc24",
  2259 => x"047c7c00",
  2260 => x"00080c04",
  2261 => x"545c4800",
  2262 => x"00207454",
  2263 => x"7f3f0400",
  2264 => x"00004444",
  2265 => x"407c3c00",
  2266 => x"007c7c40",
  2267 => x"603c1c00",
  2268 => x"001c3c60",
  2269 => x"30607c3c",
  2270 => x"003c7c60",
  2271 => x"10386c44",
  2272 => x"00446c38",
  2273 => x"e0bc1c00",
  2274 => x"001c3c60",
  2275 => x"74644400",
  2276 => x"00444c5c",
  2277 => x"3e080800",
  2278 => x"00414177",
  2279 => x"7f000000",
  2280 => x"0000007f",
  2281 => x"77414100",
  2282 => x"0008083e",
  2283 => x"03010102",
  2284 => x"00010202",
  2285 => x"7f7f7f7f",
  2286 => x"007f7f7f",
  2287 => x"1c1c0808",
  2288 => x"7f7f3e3e",
  2289 => x"3e3e7f7f",
  2290 => x"08081c1c",
  2291 => x"7c181000",
  2292 => x"0010187c",
  2293 => x"7c301000",
  2294 => x"0010307c",
  2295 => x"60603010",
  2296 => x"00061e78",
  2297 => x"183c6642",
  2298 => x"0042663c",
  2299 => x"c26a3878",
  2300 => x"00386cc6",
  2301 => x"60000060",
  2302 => x"00600000",
  2303 => x"5c5b5e0e",
  2304 => x"86fc0e5d",
  2305 => x"fbc27e71",
  2306 => x"c04cbfc8",
  2307 => x"c41ec04b",
  2308 => x"c402ab66",
  2309 => x"c24dc087",
  2310 => x"754dc187",
  2311 => x"ee49731e",
  2312 => x"86c887e1",
  2313 => x"ef49e0c0",
  2314 => x"a4c487ea",
  2315 => x"f0496a4a",
  2316 => x"c8f187f1",
  2317 => x"c184cc87",
  2318 => x"abb7c883",
  2319 => x"87cdff04",
  2320 => x"4d268efc",
  2321 => x"4b264c26",
  2322 => x"711e4f26",
  2323 => x"ccfbc24a",
  2324 => x"ccfbc25a",
  2325 => x"4978c748",
  2326 => x"2687e1fe",
  2327 => x"1e731e4f",
  2328 => x"0bfc4b71",
  2329 => x"4a730b7b",
  2330 => x"c0c19ac1",
  2331 => x"c5ed49a2",
  2332 => x"ccdfc287",
  2333 => x"264b265b",
  2334 => x"4a711e4f",
  2335 => x"721e66c4",
  2336 => x"87cbec49",
  2337 => x"4f268efc",
  2338 => x"48d4ff1e",
  2339 => x"ff78ffc3",
  2340 => x"e1c048d0",
  2341 => x"48d4ff78",
  2342 => x"487178c1",
  2343 => x"d4ff30c4",
  2344 => x"d0ff7808",
  2345 => x"78e0c048",
  2346 => x"5e0e4f26",
  2347 => x"0e5d5c5b",
  2348 => x"a6c886ec",
  2349 => x"c478c048",
  2350 => x"78bfec80",
  2351 => x"fbc280f8",
  2352 => x"c278bfc8",
  2353 => x"4cbfd0fb",
  2354 => x"c24dbfe8",
  2355 => x"49bfc8df",
  2356 => x"c787c7e4",
  2357 => x"87ffe849",
  2358 => x"99c24970",
  2359 => x"c287d005",
  2360 => x"49bfc0df",
  2361 => x"66ccb9ff",
  2362 => x"0299c199",
  2363 => x"c887cbc2",
  2364 => x"c8ff48a6",
  2365 => x"49c778bf",
  2366 => x"7087dce8",
  2367 => x"717e7449",
  2368 => x"87cd0599",
  2369 => x"c14966cc",
  2370 => x"717e7499",
  2371 => x"c4c10299",
  2372 => x"4cc8ff87",
  2373 => x"cc4b66c8",
  2374 => x"bfec48a6",
  2375 => x"87fae278",
  2376 => x"6c5ba6cc",
  2377 => x"d4887348",
  2378 => x"e8cf58a6",
  2379 => x"87d106a8",
  2380 => x"bffcdec2",
  2381 => x"c2b9c149",
  2382 => x"7159c0df",
  2383 => x"6c87c9fd",
  2384 => x"e749c74b",
  2385 => x"987087d1",
  2386 => x"87cbff05",
  2387 => x"c14966cc",
  2388 => x"c2ff0599",
  2389 => x"c24c6e87",
  2390 => x"4abfc8df",
  2391 => x"dfc2bac1",
  2392 => x"0afc5acc",
  2393 => x"9ac10a7a",
  2394 => x"49a2c0c1",
  2395 => x"c187c7e9",
  2396 => x"e2e649da",
  2397 => x"48a6c887",
  2398 => x"dfc278c1",
  2399 => x"66cc48c0",
  2400 => x"c8dfc278",
  2401 => x"c7c105bf",
  2402 => x"c0c0c887",
  2403 => x"ecdec24b",
  2404 => x"144c6e7e",
  2405 => x"87ffe549",
  2406 => x"c0029870",
  2407 => x"b57387c2",
  2408 => x"052bb7c1",
  2409 => x"7587ecff",
  2410 => x"99ffc349",
  2411 => x"49c01e71",
  2412 => x"7587c6fb",
  2413 => x"29b7c849",
  2414 => x"49c11e71",
  2415 => x"c887fafa",
  2416 => x"49fdc386",
  2417 => x"c387d0e5",
  2418 => x"cae549fa",
  2419 => x"87cec787",
  2420 => x"ffc34975",
  2421 => x"2db7c899",
  2422 => x"9d75b571",
  2423 => x"87e0c002",
  2424 => x"7ebfc8ff",
  2425 => x"dfc2496e",
  2426 => x"c289bfc4",
  2427 => x"c003a9e0",
  2428 => x"4dc087c5",
  2429 => x"c287cfc0",
  2430 => x"6e48c4df",
  2431 => x"87c6c078",
  2432 => x"48c4dfc2",
  2433 => x"497578c0",
  2434 => x"c00599c8",
  2435 => x"f5c387ce",
  2436 => x"87c3e449",
  2437 => x"99c24970",
  2438 => x"87eac002",
  2439 => x"bfccfbc2",
  2440 => x"87cac002",
  2441 => x"c288c148",
  2442 => x"c058d0fb",
  2443 => x"66c487d3",
  2444 => x"80e0c148",
  2445 => x"bf6e7e70",
  2446 => x"87c5c002",
  2447 => x"7349ff4b",
  2448 => x"48a6c80f",
  2449 => x"497578c1",
  2450 => x"c00599c4",
  2451 => x"f2c387ce",
  2452 => x"87c3e349",
  2453 => x"99c24970",
  2454 => x"87f1c002",
  2455 => x"bfccfbc2",
  2456 => x"c7486e7e",
  2457 => x"c003a8b7",
  2458 => x"486e87cb",
  2459 => x"fbc280c1",
  2460 => x"d3c058d0",
  2461 => x"4866c487",
  2462 => x"7080e0c1",
  2463 => x"02bf6e7e",
  2464 => x"4b87c5c0",
  2465 => x"0f7349fe",
  2466 => x"c148a6c8",
  2467 => x"49fdc378",
  2468 => x"7087c4e2",
  2469 => x"0299c249",
  2470 => x"c287e6c0",
  2471 => x"02bfccfb",
  2472 => x"c287c9c0",
  2473 => x"c048ccfb",
  2474 => x"87d0c078",
  2475 => x"c14a66c4",
  2476 => x"026a82e0",
  2477 => x"4b87c5c0",
  2478 => x"0f7349fd",
  2479 => x"c148a6c8",
  2480 => x"49fac378",
  2481 => x"7087d0e1",
  2482 => x"0299c249",
  2483 => x"c287edc0",
  2484 => x"48bfccfb",
  2485 => x"03a8b7c7",
  2486 => x"c287c9c0",
  2487 => x"c748ccfb",
  2488 => x"87d3c078",
  2489 => x"c14866c4",
  2490 => x"7e7080e0",
  2491 => x"c002bf6e",
  2492 => x"fc4b87c5",
  2493 => x"c80f7349",
  2494 => x"78c148a6",
  2495 => x"f0c34875",
  2496 => x"487e7098",
  2497 => x"cec00598",
  2498 => x"49dac187",
  2499 => x"7087c8e0",
  2500 => x"0299c249",
  2501 => x"6e87cac1",
  2502 => x"87cdc005",
  2503 => x"ff49dac1",
  2504 => x"7087f4df",
  2505 => x"e8c00298",
  2506 => x"49bfe887",
  2507 => x"9bffc34b",
  2508 => x"7129b7c8",
  2509 => x"e1daffb3",
  2510 => x"c3497387",
  2511 => x"997199f0",
  2512 => x"87e5ff05",
  2513 => x"ff49dac1",
  2514 => x"7087ccdf",
  2515 => x"d8ff0598",
  2516 => x"ccfbc287",
  2517 => x"cc4b49bf",
  2518 => x"8366c493",
  2519 => x"73714b6b",
  2520 => x"029c740f",
  2521 => x"6c87e9c0",
  2522 => x"87e4c002",
  2523 => x"deff496c",
  2524 => x"497087e5",
  2525 => x"c00299c1",
  2526 => x"a4c487cb",
  2527 => x"ccfbc24b",
  2528 => x"4b6b49bf",
  2529 => x"0284c80f",
  2530 => x"6c87c5c0",
  2531 => x"87dcff05",
  2532 => x"c00266c8",
  2533 => x"fbc287c8",
  2534 => x"f149bfcc",
  2535 => x"8eec87de",
  2536 => x"4c264d26",
  2537 => x"4f264b26",
  2538 => x"00000010",
  2539 => x"14111258",
  2540 => x"231c1b1d",
  2541 => x"9491595a",
  2542 => x"f4ebf2f5",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000000",
  2547 => x"5c5b5e0e",
  2548 => x"4b710e5d",
  2549 => x"d04cd4ff",
  2550 => x"78c04866",
  2551 => x"ddff49d6",
  2552 => x"ffc387f2",
  2553 => x"c3496c7c",
  2554 => x"4d7199ff",
  2555 => x"99f0c349",
  2556 => x"05a9e0c1",
  2557 => x"ffc387cb",
  2558 => x"c3486c7c",
  2559 => x"0866d098",
  2560 => x"7cffc378",
  2561 => x"c8494a6c",
  2562 => x"7cffc331",
  2563 => x"b2714a6c",
  2564 => x"31c84972",
  2565 => x"6c7cffc3",
  2566 => x"72b2714a",
  2567 => x"c331c849",
  2568 => x"4a6c7cff",
  2569 => x"d0ffb271",
  2570 => x"78e0c048",
  2571 => x"c2029b73",
  2572 => x"757b7287",
  2573 => x"264d2648",
  2574 => x"264b264c",
  2575 => x"4f261e4f",
  2576 => x"5c5b5e0e",
  2577 => x"7686f80e",
  2578 => x"49a6c81e",
  2579 => x"c487fdfd",
  2580 => x"6e4b7086",
  2581 => x"01a8c348",
  2582 => x"7387f4c2",
  2583 => x"9af0c34a",
  2584 => x"02aad0c1",
  2585 => x"e0c187c7",
  2586 => x"e2c205aa",
  2587 => x"c8497387",
  2588 => x"87c30299",
  2589 => x"7387c6ff",
  2590 => x"c29cc34c",
  2591 => x"c4c105ac",
  2592 => x"4966c487",
  2593 => x"1e7131c9",
  2594 => x"c14a66c4",
  2595 => x"fbc292cc",
  2596 => x"817249d4",
  2597 => x"87d6cdfe",
  2598 => x"daff49d8",
  2599 => x"c0c887f6",
  2600 => x"cce8c21e",
  2601 => x"ece6fd49",
  2602 => x"48d0ff87",
  2603 => x"c278e0c0",
  2604 => x"cc1ecce8",
  2605 => x"ccc14a66",
  2606 => x"d4fbc292",
  2607 => x"fe817249",
  2608 => x"cc87eccb",
  2609 => x"05acc186",
  2610 => x"c487c4c1",
  2611 => x"31c94966",
  2612 => x"66c41e71",
  2613 => x"92ccc14a",
  2614 => x"49d4fbc2",
  2615 => x"ccfe8172",
  2616 => x"e8c287cc",
  2617 => x"66c81ecc",
  2618 => x"92ccc14a",
  2619 => x"49d4fbc2",
  2620 => x"c9fe8172",
  2621 => x"49d787fa",
  2622 => x"87d8d9ff",
  2623 => x"c21ec0c8",
  2624 => x"fd49cce8",
  2625 => x"cc87ebe4",
  2626 => x"48d0ff86",
  2627 => x"f878e0c0",
  2628 => x"264c268e",
  2629 => x"1e4f264b",
  2630 => x"b7c44a71",
  2631 => x"87ce03aa",
  2632 => x"ccc14972",
  2633 => x"d4fbc291",
  2634 => x"81c8c181",
  2635 => x"4f2679c0",
  2636 => x"5c5b5e0e",
  2637 => x"86fc0e5d",
  2638 => x"d4ff4a71",
  2639 => x"d44cc04b",
  2640 => x"b7c34d66",
  2641 => x"c2c201ad",
  2642 => x"029a7287",
  2643 => x"1e87ecc0",
  2644 => x"ccc14975",
  2645 => x"d4fbc291",
  2646 => x"c8807148",
  2647 => x"66c458a6",
  2648 => x"d7c3fe49",
  2649 => x"7086c487",
  2650 => x"87d40298",
  2651 => x"c8c1496e",
  2652 => x"6e79c181",
  2653 => x"6981c849",
  2654 => x"7587c54c",
  2655 => x"87d7fe49",
  2656 => x"c848d0ff",
  2657 => x"7bdd78e1",
  2658 => x"ffc34874",
  2659 => x"747b7098",
  2660 => x"29b7c849",
  2661 => x"ffc34871",
  2662 => x"747b7098",
  2663 => x"29b7d049",
  2664 => x"ffc34871",
  2665 => x"747b7098",
  2666 => x"28b7d848",
  2667 => x"7bc07b70",
  2668 => x"7b7b7b7b",
  2669 => x"7b7b7b7b",
  2670 => x"ff7b7b7b",
  2671 => x"e0c048d0",
  2672 => x"dc1e7578",
  2673 => x"f0d6ff49",
  2674 => x"fc86c487",
  2675 => x"264d268e",
  2676 => x"264b264c",
  2677 => x"001cff4f",
  2678 => x"001cff00",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
