library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testsector is
 port (
   addr : in  std_logic_vector(12 downto 0);
   clk  : in  std_logic;
   data : out std_logic_vector(7 downto 0)
   );
end entity;

architecture prom of testsector is
  type rom is array(0 to 8191) of std_logic_vector(7 downto 0);
  signal rom_data: rom := (
     X"78", X"d8", X"a2", X"ff", X"9a", X"a9", X"80", X"85",
     X"1a", X"a9", X"bb", X"85", X"1b", X"a9", X"00", X"85",
     X"18", X"85", X"19", X"a9", X"01", X"85", X"16", X"a9",
     X"1a", X"8d", X"df", X"bf", X"20", X"8e", X"e0", X"20",
     X"24", X"e1", X"20", X"66", X"e0", X"a2", X"00", X"a0",
     X"00", X"20", X"d7", X"e0", X"a9", X"b8", X"85", X"14",
     X"a9", X"e1", X"85", X"15", X"20", X"0e", X"e1", X"a5",
     X"16", X"20", X"a5", X"e0", X"a9", X"c1", X"85", X"14",
     X"a9", X"e1", X"85", X"15", X"20", X"0e", X"e1", X"a5",
     X"17", X"20", X"a5", X"e0", X"a9", X"1f", X"20", X"c0",
     X"e0", X"20", X"43", X"e1", X"a2", X"00", X"8a", X"48",
     X"bd", X"00", X"06", X"20", X"a5", X"e0", X"68", X"aa",
     X"e8", X"d0", X"f3", X"38", X"b0", X"fe", X"a9", X"e0",
     X"85", X"14", X"a9", X"bf", X"85", X"15", X"a2", X"1c",
     X"a9", X"20", X"a0", X"27", X"91", X"14", X"88", X"10",
     X"fb", X"a5", X"14", X"38", X"e9", X"28", X"85", X"14",
     X"b0", X"02", X"c6", X"15", X"ca", X"10", X"e9", X"a2",
     X"00", X"a0", X"00", X"4c", X"d7", X"e0", X"a2", X"a8",
     X"bd", X"e8", X"e1", X"9d", X"2f", X"b5", X"ca", X"d0",
     X"f7", X"a2", X"d8", X"bd", X"90", X"e2", X"9d", X"ff",
     X"b5", X"ca", X"d0", X"f7", X"60", X"48", X"4a", X"4a",
     X"4a", X"4a", X"aa", X"bd", X"d9", X"e1", X"20", X"c0",
     X"e0", X"68", X"29", X"0f", X"aa", X"bd", X"d9", X"e1",
     X"20", X"c0", X"e0", X"a9", X"2c", X"4c", X"c0", X"e0",
     X"c9", X"1f", X"d0", X"08", X"a4", X"19", X"c8", X"a2",
     X"02", X"4c", X"d7", X"e0", X"a0", X"00", X"91", X"1a",
     X"e6", X"1a", X"d0", X"02", X"e6", X"1b", X"60", X"86",
     X"18", X"84", X"19", X"a9", X"80", X"85", X"1a", X"a9",
     X"bb", X"85", X"1b", X"a9", X"00", X"85", X"05", X"84",
     X"04", X"98", X"0a", X"0a", X"18", X"65", X"04", X"0a",
     X"26", X"05", X"0a", X"26", X"05", X"0a", X"26", X"05",
     X"18", X"65", X"1a", X"85", X"1a", X"a5", X"05", X"65",
     X"1b", X"85", X"1b", X"18", X"8a", X"65", X"1a", X"85",
     X"1a", X"90", X"02", X"e6", X"1b", X"60", X"a0", X"00",
     X"b1", X"14", X"f0", X"0f", X"84", X"1d", X"20", X"c0",
     X"e0", X"a4", X"1d", X"c8", X"d0", X"f2", X"e6", X"15",
     X"4c", X"10", X"e1", X"60", X"a9", X"0c", X"8d", X"10",
     X"03", X"20", X"33", X"e1", X"ad", X"10", X"03", X"29",
     X"10", X"d0", X"f1", X"8a", X"48", X"a2", X"05", X"ca",
     X"d0", X"fd", X"ad", X"10", X"03", X"4a", X"b0", X"fa",
     X"68", X"aa", X"60", X"a9", X"06", X"85", X"15", X"a9",
     X"00", X"85", X"14", X"a0", X"04", X"84", X"1c", X"a6",
     X"17", X"ec", X"11", X"03", X"f0", X"13", X"8e", X"13",
     X"03", X"a9", X"1f", X"8d", X"10", X"03", X"a0", X"05",
     X"88", X"d0", X"fd", X"ad", X"10", X"03", X"4a", X"b0",
     X"fa", X"a0", X"03", X"88", X"d0", X"fd", X"a5", X"16",
     X"8d", X"12", X"03", X"a9", X"04", X"8d", X"14", X"03",
     X"a9", X"80", X"8d", X"10", X"03", X"a0", X"04", X"88",
     X"d0", X"fd", X"a0", X"00", X"ad", X"10", X"03", X"4a",
     X"90", X"0e", X"ad", X"18", X"03", X"30", X"f5", X"ad",
     X"13", X"03", X"91", X"14", X"c8", X"4c", X"8a", X"e1",
     X"29", X"3e", X"f0", X"1b", X"c6", X"1c", X"d0", X"af",
     X"48", X"a2", X"02", X"a0", X"16", X"20", X"d7", X"e0",
     X"a9", X"ca", X"85", X"14", X"a9", X"e1", X"85", X"15",
     X"20", X"0e", X"e1", X"68", X"4c", X"a5", X"e0", X"60",
     X"53", X"45", X"43", X"54", X"4f", X"52", X"3a", X"20",
     X"00", X"20", X"50", X"49", X"53", X"54", X"41", X"3a",
     X"20", X"00", X"c2", X"a1", X"52", X"45", X"41", X"44",
     X"20", X"45", X"52", X"52", X"4f", X"52", X"21", X"20",
     X"00", X"30", X"31", X"32", X"33", X"34", X"35", X"36",
     X"37", X"38", X"39", X"41", X"42", X"43", X"44", X"45",
     X"46", X"4c", X"4c", X"40", X"4c", X"4c", X"48", X"50",
     X"40", X"4c", X"4c", X"4c", X"40", X"40", X"40", X"40",
     X"40", X"5e", X"46", X"46", X"46", X"46", X"5e", X"40",
     X"40", X"7c", X"70", X"70", X"70", X"70", X"7c", X"40",
     X"40", X"60", X"50", X"48", X"44", X"42", X"40", X"40",
     X"40", X"40", X"40", X"5e", X"40", X"5e", X"40", X"40",
     X"40", X"40", X"40", X"40", X"4c", X"4c", X"48", X"50",
     X"40", X"40", X"40", X"5e", X"40", X"40", X"40", X"40",
     X"40", X"40", X"40", X"40", X"40", X"4c", X"4c", X"40",
     X"40", X"42", X"44", X"48", X"50", X"60", X"40", X"40",
     X"40", X"7e", X"72", X"72", X"7a", X"7a", X"7e", X"40",
     X"40", X"4c", X"5c", X"6c", X"4c", X"4c", X"4c", X"40",
     X"40", X"7e", X"46", X"46", X"7e", X"70", X"7e", X"40",
     X"40", X"7e", X"46", X"5e", X"46", X"46", X"7e", X"40",
     X"40", X"70", X"72", X"72", X"7e", X"46", X"46", X"40",
     X"40", X"7e", X"70", X"7e", X"46", X"46", X"7c", X"40",
     X"40", X"5e", X"70", X"70", X"7e", X"72", X"7e", X"40",
     X"40", X"7e", X"46", X"4c", X"4c", X"58", X"58", X"40",
     X"40", X"7e", X"72", X"7e", X"72", X"72", X"7e", X"40",
     X"40", X"7e", X"72", X"72", X"7e", X"46", X"7e", X"40",
     X"40", X"40", X"40", X"4c", X"40", X"4c", X"40", X"40",
     X"40", X"40", X"40", X"40", X"40", X"40", X"40", X"40",
     X"40", X"7c", X"72", X"72", X"7e", X"72", X"72", X"40",
     X"40", X"7c", X"72", X"7c", X"72", X"72", X"7c", X"40",
     X"40", X"7e", X"70", X"70", X"70", X"70", X"7e", X"40",
     X"40", X"7c", X"72", X"72", X"72", X"72", X"7c", X"40",
     X"40", X"7e", X"70", X"78", X"70", X"70", X"7e", X"40",
     X"40", X"7e", X"70", X"7c", X"70", X"70", X"70", X"40",
     X"40", X"7e", X"70", X"70", X"76", X"72", X"7e", X"40",
     X"40", X"72", X"72", X"7e", X"72", X"72", X"72", X"40",
     X"40", X"7c", X"58", X"58", X"58", X"58", X"7c", X"40",
     X"40", X"5e", X"46", X"46", X"46", X"66", X"5c", X"40",
     X"40", X"72", X"74", X"78", X"74", X"72", X"72", X"40",
     X"40", X"70", X"70", X"70", X"70", X"70", X"7e", X"40",
     X"40", X"7c", X"6a", X"6a", X"62", X"72", X"72", X"40",
     X"40", X"72", X"7a", X"76", X"72", X"72", X"72", X"40",
     X"40", X"5e", X"72", X"72", X"72", X"72", X"7e", X"40",
     X"40", X"7c", X"72", X"72", X"7c", X"70", X"70", X"40",
     X"40", X"5e", X"72", X"72", X"72", X"74", X"7a", X"40",
     X"40", X"7c", X"72", X"72", X"7c", X"72", X"72", X"40",
     X"40", X"7e", X"70", X"7e", X"46", X"46", X"7e", X"40",
     X"40", X"7c", X"58", X"58", X"58", X"58", X"58", X"40",
     X"40", X"72", X"72", X"72", X"72", X"72", X"7c", X"40",
     X"40", X"72", X"72", X"72", X"72", X"74", X"78", X"40",
     X"40", X"72", X"72", X"62", X"6a", X"6a", X"7c", X"40",
     X"40", X"62", X"54", X"48", X"48", X"54", X"62", X"40",
     X"40", X"64", X"64", X"64", X"58", X"58", X"58", X"40",
     X"40", X"7e", X"46", X"4c", X"58", X"70", X"7e", X"40",
     X"40", X"e6", X"16", X"a5", X"16", X"c9", X"12", X"d0",
     X"06", X"a9", X"01", X"85", X"16", X"e6", X"17", X"68",
     X"68", X"68", X"4c", X"22", X"e0", X"40", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"69", X"e3", X"00", X"e0", X"7d", X"e3");

begin

process (clk)
  begin
    if rising_edge(clk) then
      data <= rom_data(TO_INTEGER(unsigned(addr)));
    end if;
  end process;

end architecture;
