
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"c8",x"78",x"c0",x"48"),
     1 => (x"87",x"c5",x"02",x"66"),
     2 => (x"c2",x"49",x"ff",x"c3"),
     3 => (x"c2",x"49",x"c0",x"87"),
     4 => (x"cc",x"59",x"e0",x"fb"),
     5 => (x"87",x"c6",x"02",x"66"),
     6 => (x"4a",x"d5",x"d5",x"c5"),
     7 => (x"ff",x"cf",x"87",x"c4"),
     8 => (x"fb",x"c2",x"4a",x"ff"),
     9 => (x"fb",x"c2",x"5a",x"e4"),
    10 => (x"78",x"c1",x"48",x"e4"),
    11 => (x"4f",x"26",x"4b",x"26"),
    12 => (x"5c",x"5b",x"5e",x"0e"),
    13 => (x"4d",x"71",x"0e",x"5d"),
    14 => (x"bf",x"e0",x"fb",x"c2"),
    15 => (x"02",x"9d",x"75",x"4b"),
    16 => (x"c8",x"49",x"87",x"cb"),
    17 => (x"d8",x"ff",x"c1",x"91"),
    18 => (x"c4",x"82",x"71",x"4a"),
    19 => (x"d8",x"c3",x"c2",x"87"),
    20 => (x"12",x"4c",x"c0",x"4a"),
    21 => (x"c2",x"99",x"73",x"49"),
    22 => (x"48",x"bf",x"dc",x"fb"),
    23 => (x"d4",x"ff",x"b8",x"71"),
    24 => (x"b7",x"c1",x"78",x"08"),
    25 => (x"b7",x"c8",x"84",x"2b"),
    26 => (x"87",x"e7",x"04",x"ac"),
    27 => (x"bf",x"d8",x"fb",x"c2"),
    28 => (x"c2",x"80",x"c8",x"48"),
    29 => (x"26",x"58",x"dc",x"fb"),
    30 => (x"26",x"4c",x"26",x"4d"),
    31 => (x"1e",x"4f",x"26",x"4b"),
    32 => (x"4b",x"71",x"1e",x"73"),
    33 => (x"02",x"9a",x"4a",x"13"),
    34 => (x"49",x"72",x"87",x"cb"),
    35 => (x"13",x"87",x"e1",x"fe"),
    36 => (x"f5",x"05",x"9a",x"4a"),
    37 => (x"26",x"4b",x"26",x"87"),
    38 => (x"fb",x"c2",x"1e",x"4f"),
    39 => (x"c2",x"49",x"bf",x"d8"),
    40 => (x"c1",x"48",x"d8",x"fb"),
    41 => (x"c0",x"c4",x"78",x"a1"),
    42 => (x"db",x"03",x"a9",x"b7"),
    43 => (x"48",x"d4",x"ff",x"87"),
    44 => (x"bf",x"dc",x"fb",x"c2"),
    45 => (x"d8",x"fb",x"c2",x"78"),
    46 => (x"fb",x"c2",x"49",x"bf"),
    47 => (x"a1",x"c1",x"48",x"d8"),
    48 => (x"b7",x"c0",x"c4",x"78"),
    49 => (x"87",x"e5",x"04",x"a9"),
    50 => (x"c8",x"48",x"d0",x"ff"),
    51 => (x"e4",x"fb",x"c2",x"78"),
    52 => (x"26",x"78",x"c0",x"48"),
    53 => (x"00",x"00",x"00",x"4f"),
    54 => (x"00",x"00",x"00",x"00"),
    55 => (x"00",x"00",x"00",x"00"),
    56 => (x"5f",x"00",x"00",x"00"),
    57 => (x"00",x"00",x"00",x"5f"),
    58 => (x"00",x"03",x"03",x"00"),
    59 => (x"00",x"00",x"03",x"03"),
    60 => (x"14",x"7f",x"7f",x"14"),
    61 => (x"00",x"14",x"7f",x"7f"),
    62 => (x"6b",x"2e",x"24",x"00"),
    63 => (x"00",x"12",x"3a",x"6b"),
    64 => (x"18",x"36",x"6a",x"4c"),
    65 => (x"00",x"32",x"56",x"6c"),
    66 => (x"59",x"4f",x"7e",x"30"),
    67 => (x"40",x"68",x"3a",x"77"),
    68 => (x"07",x"04",x"00",x"00"),
    69 => (x"00",x"00",x"00",x"03"),
    70 => (x"3e",x"1c",x"00",x"00"),
    71 => (x"00",x"00",x"41",x"63"),
    72 => (x"63",x"41",x"00",x"00"),
    73 => (x"00",x"00",x"1c",x"3e"),
    74 => (x"1c",x"3e",x"2a",x"08"),
    75 => (x"08",x"2a",x"3e",x"1c"),
    76 => (x"3e",x"08",x"08",x"00"),
    77 => (x"00",x"08",x"08",x"3e"),
    78 => (x"e0",x"80",x"00",x"00"),
    79 => (x"00",x"00",x"00",x"60"),
    80 => (x"08",x"08",x"08",x"00"),
    81 => (x"00",x"08",x"08",x"08"),
    82 => (x"60",x"00",x"00",x"00"),
    83 => (x"00",x"00",x"00",x"60"),
    84 => (x"18",x"30",x"60",x"40"),
    85 => (x"01",x"03",x"06",x"0c"),
    86 => (x"59",x"7f",x"3e",x"00"),
    87 => (x"00",x"3e",x"7f",x"4d"),
    88 => (x"7f",x"06",x"04",x"00"),
    89 => (x"00",x"00",x"00",x"7f"),
    90 => (x"71",x"63",x"42",x"00"),
    91 => (x"00",x"46",x"4f",x"59"),
    92 => (x"49",x"63",x"22",x"00"),
    93 => (x"00",x"36",x"7f",x"49"),
    94 => (x"13",x"16",x"1c",x"18"),
    95 => (x"00",x"10",x"7f",x"7f"),
    96 => (x"45",x"67",x"27",x"00"),
    97 => (x"00",x"39",x"7d",x"45"),
    98 => (x"4b",x"7e",x"3c",x"00"),
    99 => (x"00",x"30",x"79",x"49"),
   100 => (x"71",x"01",x"01",x"00"),
   101 => (x"00",x"07",x"0f",x"79"),
   102 => (x"49",x"7f",x"36",x"00"),
   103 => (x"00",x"36",x"7f",x"49"),
   104 => (x"49",x"4f",x"06",x"00"),
   105 => (x"00",x"1e",x"3f",x"69"),
   106 => (x"66",x"00",x"00",x"00"),
   107 => (x"00",x"00",x"00",x"66"),
   108 => (x"e6",x"80",x"00",x"00"),
   109 => (x"00",x"00",x"00",x"66"),
   110 => (x"14",x"08",x"08",x"00"),
   111 => (x"00",x"22",x"22",x"14"),
   112 => (x"14",x"14",x"14",x"00"),
   113 => (x"00",x"14",x"14",x"14"),
   114 => (x"14",x"22",x"22",x"00"),
   115 => (x"00",x"08",x"08",x"14"),
   116 => (x"51",x"03",x"02",x"00"),
   117 => (x"00",x"06",x"0f",x"59"),
   118 => (x"5d",x"41",x"7f",x"3e"),
   119 => (x"00",x"1e",x"1f",x"55"),
   120 => (x"09",x"7f",x"7e",x"00"),
   121 => (x"00",x"7e",x"7f",x"09"),
   122 => (x"49",x"7f",x"7f",x"00"),
   123 => (x"00",x"36",x"7f",x"49"),
   124 => (x"63",x"3e",x"1c",x"00"),
   125 => (x"00",x"41",x"41",x"41"),
   126 => (x"41",x"7f",x"7f",x"00"),
   127 => (x"00",x"1c",x"3e",x"63"),
   128 => (x"49",x"7f",x"7f",x"00"),
   129 => (x"00",x"41",x"41",x"49"),
   130 => (x"09",x"7f",x"7f",x"00"),
   131 => (x"00",x"01",x"01",x"09"),
   132 => (x"41",x"7f",x"3e",x"00"),
   133 => (x"00",x"7a",x"7b",x"49"),
   134 => (x"08",x"7f",x"7f",x"00"),
   135 => (x"00",x"7f",x"7f",x"08"),
   136 => (x"7f",x"41",x"00",x"00"),
   137 => (x"00",x"00",x"41",x"7f"),
   138 => (x"40",x"60",x"20",x"00"),
   139 => (x"00",x"3f",x"7f",x"40"),
   140 => (x"1c",x"08",x"7f",x"7f"),
   141 => (x"00",x"41",x"63",x"36"),
   142 => (x"40",x"7f",x"7f",x"00"),
   143 => (x"00",x"40",x"40",x"40"),
   144 => (x"0c",x"06",x"7f",x"7f"),
   145 => (x"00",x"7f",x"7f",x"06"),
   146 => (x"0c",x"06",x"7f",x"7f"),
   147 => (x"00",x"7f",x"7f",x"18"),
   148 => (x"41",x"7f",x"3e",x"00"),
   149 => (x"00",x"3e",x"7f",x"41"),
   150 => (x"09",x"7f",x"7f",x"00"),
   151 => (x"00",x"06",x"0f",x"09"),
   152 => (x"61",x"41",x"7f",x"3e"),
   153 => (x"00",x"40",x"7e",x"7f"),
   154 => (x"09",x"7f",x"7f",x"00"),
   155 => (x"00",x"66",x"7f",x"19"),
   156 => (x"4d",x"6f",x"26",x"00"),
   157 => (x"00",x"32",x"7b",x"59"),
   158 => (x"7f",x"01",x"01",x"00"),
   159 => (x"00",x"01",x"01",x"7f"),
   160 => (x"40",x"7f",x"3f",x"00"),
   161 => (x"00",x"3f",x"7f",x"40"),
   162 => (x"70",x"3f",x"0f",x"00"),
   163 => (x"00",x"0f",x"3f",x"70"),
   164 => (x"18",x"30",x"7f",x"7f"),
   165 => (x"00",x"7f",x"7f",x"30"),
   166 => (x"1c",x"36",x"63",x"41"),
   167 => (x"41",x"63",x"36",x"1c"),
   168 => (x"7c",x"06",x"03",x"01"),
   169 => (x"01",x"03",x"06",x"7c"),
   170 => (x"4d",x"59",x"71",x"61"),
   171 => (x"00",x"41",x"43",x"47"),
   172 => (x"7f",x"7f",x"00",x"00"),
   173 => (x"00",x"00",x"41",x"41"),
   174 => (x"0c",x"06",x"03",x"01"),
   175 => (x"40",x"60",x"30",x"18"),
   176 => (x"41",x"41",x"00",x"00"),
   177 => (x"00",x"00",x"7f",x"7f"),
   178 => (x"03",x"06",x"0c",x"08"),
   179 => (x"00",x"08",x"0c",x"06"),
   180 => (x"80",x"80",x"80",x"80"),
   181 => (x"00",x"80",x"80",x"80"),
   182 => (x"03",x"00",x"00",x"00"),
   183 => (x"00",x"00",x"04",x"07"),
   184 => (x"54",x"74",x"20",x"00"),
   185 => (x"00",x"78",x"7c",x"54"),
   186 => (x"44",x"7f",x"7f",x"00"),
   187 => (x"00",x"38",x"7c",x"44"),
   188 => (x"44",x"7c",x"38",x"00"),
   189 => (x"00",x"00",x"44",x"44"),
   190 => (x"44",x"7c",x"38",x"00"),
   191 => (x"00",x"7f",x"7f",x"44"),
   192 => (x"54",x"7c",x"38",x"00"),
   193 => (x"00",x"18",x"5c",x"54"),
   194 => (x"7f",x"7e",x"04",x"00"),
   195 => (x"00",x"00",x"05",x"05"),
   196 => (x"a4",x"bc",x"18",x"00"),
   197 => (x"00",x"7c",x"fc",x"a4"),
   198 => (x"04",x"7f",x"7f",x"00"),
   199 => (x"00",x"78",x"7c",x"04"),
   200 => (x"3d",x"00",x"00",x"00"),
   201 => (x"00",x"00",x"40",x"7d"),
   202 => (x"80",x"80",x"80",x"00"),
   203 => (x"00",x"00",x"7d",x"fd"),
   204 => (x"10",x"7f",x"7f",x"00"),
   205 => (x"00",x"44",x"6c",x"38"),
   206 => (x"3f",x"00",x"00",x"00"),
   207 => (x"00",x"00",x"40",x"7f"),
   208 => (x"18",x"0c",x"7c",x"7c"),
   209 => (x"00",x"78",x"7c",x"0c"),
   210 => (x"04",x"7c",x"7c",x"00"),
   211 => (x"00",x"78",x"7c",x"04"),
   212 => (x"44",x"7c",x"38",x"00"),
   213 => (x"00",x"38",x"7c",x"44"),
   214 => (x"24",x"fc",x"fc",x"00"),
   215 => (x"00",x"18",x"3c",x"24"),
   216 => (x"24",x"3c",x"18",x"00"),
   217 => (x"00",x"fc",x"fc",x"24"),
   218 => (x"04",x"7c",x"7c",x"00"),
   219 => (x"00",x"08",x"0c",x"04"),
   220 => (x"54",x"5c",x"48",x"00"),
   221 => (x"00",x"20",x"74",x"54"),
   222 => (x"7f",x"3f",x"04",x"00"),
   223 => (x"00",x"00",x"44",x"44"),
   224 => (x"40",x"7c",x"3c",x"00"),
   225 => (x"00",x"7c",x"7c",x"40"),
   226 => (x"60",x"3c",x"1c",x"00"),
   227 => (x"00",x"1c",x"3c",x"60"),
   228 => (x"30",x"60",x"7c",x"3c"),
   229 => (x"00",x"3c",x"7c",x"60"),
   230 => (x"10",x"38",x"6c",x"44"),
   231 => (x"00",x"44",x"6c",x"38"),
   232 => (x"e0",x"bc",x"1c",x"00"),
   233 => (x"00",x"1c",x"3c",x"60"),
   234 => (x"74",x"64",x"44",x"00"),
   235 => (x"00",x"44",x"4c",x"5c"),
   236 => (x"3e",x"08",x"08",x"00"),
   237 => (x"00",x"41",x"41",x"77"),
   238 => (x"7f",x"00",x"00",x"00"),
   239 => (x"00",x"00",x"00",x"7f"),
   240 => (x"77",x"41",x"41",x"00"),
   241 => (x"00",x"08",x"08",x"3e"),
   242 => (x"03",x"01",x"01",x"02"),
   243 => (x"00",x"01",x"02",x"02"),
   244 => (x"7f",x"7f",x"7f",x"7f"),
   245 => (x"00",x"7f",x"7f",x"7f"),
   246 => (x"1c",x"1c",x"08",x"08"),
   247 => (x"7f",x"7f",x"3e",x"3e"),
   248 => (x"3e",x"3e",x"7f",x"7f"),
   249 => (x"08",x"08",x"1c",x"1c"),
   250 => (x"7c",x"18",x"10",x"00"),
   251 => (x"00",x"10",x"18",x"7c"),
   252 => (x"7c",x"30",x"10",x"00"),
   253 => (x"00",x"10",x"30",x"7c"),
   254 => (x"60",x"60",x"30",x"10"),
   255 => (x"00",x"06",x"1e",x"78"),
   256 => (x"18",x"3c",x"66",x"42"),
   257 => (x"00",x"42",x"66",x"3c"),
   258 => (x"c2",x"6a",x"38",x"78"),
   259 => (x"00",x"38",x"6c",x"c6"),
   260 => (x"60",x"00",x"00",x"60"),
   261 => (x"00",x"60",x"00",x"00"),
   262 => (x"5c",x"5b",x"5e",x"0e"),
   263 => (x"86",x"fc",x"0e",x"5d"),
   264 => (x"c2",x"59",x"a6",x"c4"),
   265 => (x"4c",x"bf",x"ec",x"fb"),
   266 => (x"1e",x"c0",x"4b",x"c0"),
   267 => (x"02",x"ab",x"66",x"c4"),
   268 => (x"4d",x"c0",x"87",x"c4"),
   269 => (x"4d",x"c1",x"87",x"c2"),
   270 => (x"49",x"73",x"1e",x"75"),
   271 => (x"c8",x"87",x"e0",x"ee"),
   272 => (x"49",x"e0",x"c0",x"86"),
   273 => (x"c4",x"87",x"e9",x"ef"),
   274 => (x"49",x"6a",x"4a",x"a4"),
   275 => (x"f1",x"87",x"f0",x"f0"),
   276 => (x"84",x"cc",x"87",x"c7"),
   277 => (x"b7",x"c8",x"83",x"c1"),
   278 => (x"cd",x"ff",x"04",x"ab"),
   279 => (x"26",x"8e",x"fc",x"87"),
   280 => (x"26",x"4c",x"26",x"4d"),
   281 => (x"1e",x"4f",x"26",x"4b"),
   282 => (x"fb",x"c2",x"4a",x"71"),
   283 => (x"fb",x"c2",x"5a",x"f0"),
   284 => (x"78",x"c7",x"48",x"f0"),
   285 => (x"87",x"e0",x"fe",x"49"),
   286 => (x"73",x"1e",x"4f",x"26"),
   287 => (x"fc",x"4b",x"71",x"1e"),
   288 => (x"73",x"0b",x"7b",x"0b"),
   289 => (x"c1",x"9a",x"c1",x"4a"),
   290 => (x"ed",x"49",x"a2",x"c0"),
   291 => (x"df",x"c2",x"87",x"c4"),
   292 => (x"4b",x"26",x"5b",x"f0"),
   293 => (x"71",x"1e",x"4f",x"26"),
   294 => (x"1e",x"66",x"c4",x"4a"),
   295 => (x"ca",x"ec",x"49",x"72"),
   296 => (x"26",x"8e",x"fc",x"87"),
   297 => (x"d4",x"ff",x"1e",x"4f"),
   298 => (x"78",x"ff",x"c3",x"48"),
   299 => (x"c0",x"48",x"d0",x"ff"),
   300 => (x"d4",x"ff",x"78",x"e1"),
   301 => (x"71",x"78",x"c1",x"48"),
   302 => (x"ff",x"30",x"c4",x"48"),
   303 => (x"ff",x"78",x"08",x"d4"),
   304 => (x"e0",x"c0",x"48",x"d0"),
   305 => (x"0e",x"4f",x"26",x"78"),
   306 => (x"5d",x"5c",x"5b",x"5e"),
   307 => (x"c8",x"86",x"ec",x"0e"),
   308 => (x"78",x"c0",x"48",x"a6"),
   309 => (x"bf",x"ec",x"80",x"c4"),
   310 => (x"c2",x"80",x"f8",x"78"),
   311 => (x"78",x"bf",x"ec",x"fb"),
   312 => (x"bf",x"f4",x"fb",x"c2"),
   313 => (x"4d",x"bf",x"e8",x"4c"),
   314 => (x"bf",x"ec",x"df",x"c2"),
   315 => (x"87",x"c5",x"e4",x"49"),
   316 => (x"fe",x"e8",x"49",x"c7"),
   317 => (x"c2",x"49",x"70",x"87"),
   318 => (x"87",x"d0",x"05",x"99"),
   319 => (x"bf",x"e4",x"df",x"c2"),
   320 => (x"cc",x"b9",x"ff",x"49"),
   321 => (x"99",x"c1",x"99",x"66"),
   322 => (x"87",x"cd",x"c2",x"02"),
   323 => (x"ff",x"48",x"a6",x"c8"),
   324 => (x"c7",x"78",x"bf",x"c8"),
   325 => (x"87",x"db",x"e8",x"49"),
   326 => (x"a6",x"c4",x"49",x"70"),
   327 => (x"05",x"99",x"71",x"5c"),
   328 => (x"66",x"cc",x"87",x"ce"),
   329 => (x"c4",x"99",x"c1",x"49"),
   330 => (x"99",x"71",x"5c",x"a6"),
   331 => (x"87",x"c4",x"c1",x"02"),
   332 => (x"c8",x"4c",x"c8",x"ff"),
   333 => (x"a6",x"cc",x"4b",x"66"),
   334 => (x"78",x"bf",x"ec",x"48"),
   335 => (x"cc",x"87",x"f6",x"e2"),
   336 => (x"48",x"6c",x"5b",x"a6"),
   337 => (x"a6",x"d4",x"88",x"73"),
   338 => (x"a8",x"e8",x"cf",x"58"),
   339 => (x"c2",x"87",x"d1",x"06"),
   340 => (x"49",x"bf",x"e0",x"df"),
   341 => (x"df",x"c2",x"b9",x"c1"),
   342 => (x"fd",x"71",x"59",x"e4"),
   343 => (x"4b",x"6c",x"87",x"c7"),
   344 => (x"ce",x"e7",x"49",x"c7"),
   345 => (x"05",x"98",x"70",x"87"),
   346 => (x"cc",x"87",x"cb",x"ff"),
   347 => (x"99",x"c1",x"49",x"66"),
   348 => (x"87",x"c2",x"ff",x"05"),
   349 => (x"df",x"c2",x"4c",x"6e"),
   350 => (x"c1",x"4a",x"bf",x"ec"),
   351 => (x"f0",x"df",x"c2",x"ba"),
   352 => (x"7a",x"0a",x"fc",x"5a"),
   353 => (x"c1",x"9a",x"c1",x"0a"),
   354 => (x"e9",x"49",x"a2",x"c0"),
   355 => (x"da",x"c1",x"87",x"c4"),
   356 => (x"87",x"df",x"e6",x"49"),
   357 => (x"c1",x"48",x"a6",x"c8"),
   358 => (x"e4",x"df",x"c2",x"78"),
   359 => (x"78",x"66",x"cc",x"48"),
   360 => (x"bf",x"ec",x"df",x"c2"),
   361 => (x"87",x"c7",x"c1",x"05"),
   362 => (x"4b",x"c0",x"c0",x"c8"),
   363 => (x"7e",x"d0",x"df",x"c2"),
   364 => (x"49",x"14",x"4c",x"6e"),
   365 => (x"70",x"87",x"fc",x"e5"),
   366 => (x"c2",x"c0",x"02",x"98"),
   367 => (x"c1",x"b5",x"73",x"87"),
   368 => (x"ff",x"05",x"2b",x"b7"),
   369 => (x"49",x"75",x"87",x"ec"),
   370 => (x"71",x"99",x"ff",x"c3"),
   371 => (x"fb",x"49",x"c0",x"1e"),
   372 => (x"49",x"75",x"87",x"c4"),
   373 => (x"71",x"29",x"b7",x"c8"),
   374 => (x"fa",x"49",x"c1",x"1e"),
   375 => (x"86",x"c8",x"87",x"f8"),
   376 => (x"e5",x"49",x"fd",x"c3"),
   377 => (x"fa",x"c3",x"87",x"cd"),
   378 => (x"87",x"c7",x"e5",x"49"),
   379 => (x"75",x"87",x"d2",x"c7"),
   380 => (x"99",x"ff",x"c3",x"49"),
   381 => (x"71",x"2d",x"b7",x"c8"),
   382 => (x"02",x"9d",x"75",x"b5"),
   383 => (x"ff",x"87",x"e0",x"c0"),
   384 => (x"6e",x"7e",x"bf",x"c8"),
   385 => (x"e8",x"df",x"c2",x"49"),
   386 => (x"e0",x"c2",x"89",x"bf"),
   387 => (x"c5",x"c0",x"03",x"a9"),
   388 => (x"c0",x"4d",x"c0",x"87"),
   389 => (x"df",x"c2",x"87",x"cf"),
   390 => (x"78",x"6e",x"48",x"e8"),
   391 => (x"c2",x"87",x"c6",x"c0"),
   392 => (x"c0",x"48",x"e8",x"df"),
   393 => (x"c8",x"49",x"75",x"78"),
   394 => (x"ce",x"c0",x"05",x"99"),
   395 => (x"49",x"f5",x"c3",x"87"),
   396 => (x"70",x"87",x"c0",x"e4"),
   397 => (x"02",x"99",x"c2",x"49"),
   398 => (x"c2",x"87",x"eb",x"c0"),
   399 => (x"02",x"bf",x"f0",x"fb"),
   400 => (x"48",x"87",x"ca",x"c0"),
   401 => (x"fb",x"c2",x"88",x"c1"),
   402 => (x"d4",x"c0",x"58",x"f4"),
   403 => (x"48",x"66",x"c4",x"87"),
   404 => (x"c4",x"80",x"e0",x"c1"),
   405 => (x"bf",x"6e",x"58",x"a6"),
   406 => (x"87",x"c5",x"c0",x"02"),
   407 => (x"73",x"49",x"ff",x"4b"),
   408 => (x"48",x"a6",x"c8",x"0f"),
   409 => (x"49",x"75",x"78",x"c1"),
   410 => (x"c0",x"05",x"99",x"c4"),
   411 => (x"f2",x"c3",x"87",x"ce"),
   412 => (x"87",x"ff",x"e2",x"49"),
   413 => (x"99",x"c2",x"49",x"70"),
   414 => (x"87",x"f2",x"c0",x"02"),
   415 => (x"bf",x"f0",x"fb",x"c2"),
   416 => (x"c7",x"48",x"6e",x"7e"),
   417 => (x"c0",x"03",x"a8",x"b7"),
   418 => (x"48",x"6e",x"87",x"cb"),
   419 => (x"fb",x"c2",x"80",x"c1"),
   420 => (x"d4",x"c0",x"58",x"f4"),
   421 => (x"48",x"66",x"c4",x"87"),
   422 => (x"c4",x"80",x"e0",x"c1"),
   423 => (x"bf",x"6e",x"58",x"a6"),
   424 => (x"87",x"c5",x"c0",x"02"),
   425 => (x"73",x"49",x"fe",x"4b"),
   426 => (x"48",x"a6",x"c8",x"0f"),
   427 => (x"fd",x"c3",x"78",x"c1"),
   428 => (x"87",x"ff",x"e1",x"49"),
   429 => (x"99",x"c2",x"49",x"70"),
   430 => (x"87",x"e6",x"c0",x"02"),
   431 => (x"bf",x"f0",x"fb",x"c2"),
   432 => (x"87",x"c9",x"c0",x"02"),
   433 => (x"48",x"f0",x"fb",x"c2"),
   434 => (x"d0",x"c0",x"78",x"c0"),
   435 => (x"4a",x"66",x"c4",x"87"),
   436 => (x"6a",x"82",x"e0",x"c1"),
   437 => (x"87",x"c5",x"c0",x"02"),
   438 => (x"73",x"49",x"fd",x"4b"),
   439 => (x"48",x"a6",x"c8",x"0f"),
   440 => (x"fa",x"c3",x"78",x"c1"),
   441 => (x"87",x"cb",x"e1",x"49"),
   442 => (x"99",x"c2",x"49",x"70"),
   443 => (x"87",x"ee",x"c0",x"02"),
   444 => (x"bf",x"f0",x"fb",x"c2"),
   445 => (x"a8",x"b7",x"c7",x"48"),
   446 => (x"87",x"c9",x"c0",x"03"),
   447 => (x"48",x"f0",x"fb",x"c2"),
   448 => (x"d4",x"c0",x"78",x"c7"),
   449 => (x"48",x"66",x"c4",x"87"),
   450 => (x"c4",x"80",x"e0",x"c1"),
   451 => (x"bf",x"6e",x"58",x"a6"),
   452 => (x"87",x"c5",x"c0",x"02"),
   453 => (x"73",x"49",x"fc",x"4b"),
   454 => (x"48",x"a6",x"c8",x"0f"),
   455 => (x"48",x"75",x"78",x"c1"),
   456 => (x"c4",x"98",x"f0",x"c3"),
   457 => (x"98",x"70",x"58",x"a6"),
   458 => (x"87",x"ce",x"c0",x"05"),
   459 => (x"e0",x"49",x"da",x"c1"),
   460 => (x"49",x"70",x"87",x"c1"),
   461 => (x"c1",x"02",x"99",x"c2"),
   462 => (x"05",x"6e",x"87",x"ca"),
   463 => (x"c1",x"87",x"cd",x"c0"),
   464 => (x"df",x"ff",x"49",x"da"),
   465 => (x"98",x"70",x"87",x"ed"),
   466 => (x"87",x"e8",x"c0",x"02"),
   467 => (x"4b",x"49",x"bf",x"e8"),
   468 => (x"c8",x"9b",x"ff",x"c3"),
   469 => (x"b3",x"71",x"29",x"b7"),
   470 => (x"87",x"d9",x"da",x"ff"),
   471 => (x"f0",x"c3",x"49",x"73"),
   472 => (x"05",x"99",x"71",x"99"),
   473 => (x"c1",x"87",x"e5",x"ff"),
   474 => (x"df",x"ff",x"49",x"da"),
   475 => (x"98",x"70",x"87",x"c5"),
   476 => (x"87",x"d8",x"ff",x"05"),
   477 => (x"bf",x"f0",x"fb",x"c2"),
   478 => (x"93",x"cc",x"4b",x"49"),
   479 => (x"6b",x"83",x"66",x"c4"),
   480 => (x"0f",x"73",x"71",x"4b"),
   481 => (x"c0",x"02",x"9c",x"74"),
   482 => (x"02",x"6c",x"87",x"e9"),
   483 => (x"6c",x"87",x"e4",x"c0"),
   484 => (x"de",x"de",x"ff",x"49"),
   485 => (x"c1",x"49",x"70",x"87"),
   486 => (x"cb",x"c0",x"02",x"99"),
   487 => (x"4b",x"a4",x"c4",x"87"),
   488 => (x"bf",x"f0",x"fb",x"c2"),
   489 => (x"0f",x"4b",x"6b",x"49"),
   490 => (x"c0",x"02",x"84",x"c8"),
   491 => (x"05",x"6c",x"87",x"c5"),
   492 => (x"c8",x"87",x"dc",x"ff"),
   493 => (x"c8",x"c0",x"02",x"66"),
   494 => (x"f0",x"fb",x"c2",x"87"),
   495 => (x"d7",x"f1",x"49",x"bf"),
   496 => (x"26",x"8e",x"ec",x"87"),
   497 => (x"26",x"4c",x"26",x"4d"),
   498 => (x"00",x"4f",x"26",x"4b"),
   499 => (x"00",x"00",x"00",x"10"),
   500 => (x"14",x"11",x"12",x"58"),
   501 => (x"23",x"1c",x"1b",x"1d"),
   502 => (x"94",x"91",x"59",x"5a"),
   503 => (x"f4",x"eb",x"f2",x"f5"),
   504 => (x"00",x"00",x"00",x"00"),
   505 => (x"00",x"00",x"00",x"00"),
   506 => (x"00",x"00",x"00",x"00"),
   507 => (x"00",x"00",x"00",x"00"),
   508 => (x"5c",x"5b",x"5e",x"0e"),
   509 => (x"4b",x"71",x"0e",x"5d"),
   510 => (x"d0",x"4c",x"d4",x"ff"),
   511 => (x"78",x"c0",x"48",x"66"),
   512 => (x"dd",x"ff",x"49",x"d6"),
   513 => (x"ff",x"c3",x"87",x"ea"),
   514 => (x"c3",x"49",x"6c",x"7c"),
   515 => (x"4d",x"71",x"99",x"ff"),
   516 => (x"99",x"f0",x"c3",x"49"),
   517 => (x"05",x"a9",x"e0",x"c1"),
   518 => (x"ff",x"c3",x"87",x"cb"),
   519 => (x"c3",x"48",x"6c",x"7c"),
   520 => (x"08",x"66",x"d0",x"98"),
   521 => (x"7c",x"ff",x"c3",x"78"),
   522 => (x"c8",x"49",x"4a",x"6c"),
   523 => (x"7c",x"ff",x"c3",x"31"),
   524 => (x"b2",x"71",x"4a",x"6c"),
   525 => (x"31",x"c8",x"49",x"72"),
   526 => (x"6c",x"7c",x"ff",x"c3"),
   527 => (x"72",x"b2",x"71",x"4a"),
   528 => (x"c3",x"31",x"c8",x"49"),
   529 => (x"4a",x"6c",x"7c",x"ff"),
   530 => (x"d0",x"ff",x"b2",x"71"),
   531 => (x"78",x"e0",x"c0",x"48"),
   532 => (x"c2",x"02",x"9b",x"73"),
   533 => (x"75",x"7b",x"72",x"87"),
   534 => (x"26",x"4d",x"26",x"48"),
   535 => (x"26",x"4b",x"26",x"4c"),
   536 => (x"4f",x"26",x"1e",x"4f"),
   537 => (x"5c",x"5b",x"5e",x"0e"),
   538 => (x"76",x"86",x"f8",x"0e"),
   539 => (x"80",x"c4",x"48",x"1e"),
   540 => (x"fb",x"fd",x"49",x"70"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"c3",x"48",x"6e",x"4b"),
   543 => (x"f4",x"c2",x"01",x"a8"),
   544 => (x"c3",x"4a",x"73",x"87"),
   545 => (x"d0",x"c1",x"9a",x"f0"),
   546 => (x"87",x"c7",x"02",x"aa"),
   547 => (x"05",x"aa",x"e0",x"c1"),
   548 => (x"73",x"87",x"e2",x"c2"),
   549 => (x"02",x"99",x"c8",x"49"),
   550 => (x"c4",x"ff",x"87",x"c3"),
   551 => (x"c3",x"4c",x"73",x"87"),
   552 => (x"05",x"ac",x"c2",x"9c"),
   553 => (x"c4",x"87",x"c4",x"c1"),
   554 => (x"31",x"c9",x"49",x"66"),
   555 => (x"66",x"c4",x"1e",x"71"),
   556 => (x"92",x"cc",x"c1",x"4a"),
   557 => (x"49",x"f8",x"fb",x"c2"),
   558 => (x"cc",x"fe",x"81",x"72"),
   559 => (x"49",x"d8",x"87",x"fe"),
   560 => (x"87",x"ec",x"da",x"ff"),
   561 => (x"c2",x"1e",x"c0",x"c8"),
   562 => (x"fd",x"49",x"f0",x"e8"),
   563 => (x"ff",x"87",x"d0",x"e6"),
   564 => (x"e0",x"c0",x"48",x"d0"),
   565 => (x"f0",x"e8",x"c2",x"78"),
   566 => (x"4a",x"66",x"cc",x"1e"),
   567 => (x"c2",x"92",x"cc",x"c1"),
   568 => (x"72",x"49",x"f8",x"fb"),
   569 => (x"d4",x"cb",x"fe",x"81"),
   570 => (x"c1",x"86",x"cc",x"87"),
   571 => (x"c4",x"c1",x"05",x"ac"),
   572 => (x"49",x"66",x"c4",x"87"),
   573 => (x"1e",x"71",x"31",x"c9"),
   574 => (x"c1",x"4a",x"66",x"c4"),
   575 => (x"fb",x"c2",x"92",x"cc"),
   576 => (x"81",x"72",x"49",x"f8"),
   577 => (x"87",x"f4",x"cb",x"fe"),
   578 => (x"1e",x"f0",x"e8",x"c2"),
   579 => (x"c1",x"4a",x"66",x"c8"),
   580 => (x"fb",x"c2",x"92",x"cc"),
   581 => (x"81",x"72",x"49",x"f8"),
   582 => (x"87",x"e2",x"c9",x"fe"),
   583 => (x"d9",x"ff",x"49",x"d7"),
   584 => (x"c0",x"c8",x"87",x"ce"),
   585 => (x"f0",x"e8",x"c2",x"1e"),
   586 => (x"cf",x"e4",x"fd",x"49"),
   587 => (x"ff",x"86",x"cc",x"87"),
   588 => (x"e0",x"c0",x"48",x"d0"),
   589 => (x"26",x"8e",x"f8",x"78"),
   590 => (x"26",x"4b",x"26",x"4c"),
   591 => (x"4a",x"71",x"1e",x"4f"),
   592 => (x"03",x"aa",x"b7",x"c4"),
   593 => (x"49",x"72",x"87",x"ce"),
   594 => (x"c2",x"91",x"cc",x"c1"),
   595 => (x"c1",x"81",x"f8",x"fb"),
   596 => (x"79",x"c0",x"81",x"c8"),
   597 => (x"5e",x"0e",x"4f",x"26"),
   598 => (x"0e",x"5d",x"5c",x"5b"),
   599 => (x"4a",x"71",x"86",x"fc"),
   600 => (x"c0",x"4b",x"d4",x"ff"),
   601 => (x"4d",x"66",x"d4",x"4c"),
   602 => (x"01",x"ad",x"b7",x"c3"),
   603 => (x"72",x"87",x"c2",x"c2"),
   604 => (x"ec",x"c0",x"02",x"9a"),
   605 => (x"49",x"75",x"1e",x"87"),
   606 => (x"c2",x"91",x"cc",x"c1"),
   607 => (x"71",x"48",x"f8",x"fb"),
   608 => (x"58",x"a6",x"c8",x"80"),
   609 => (x"fe",x"49",x"66",x"c4"),
   610 => (x"c4",x"87",x"fd",x"c2"),
   611 => (x"02",x"98",x"70",x"86"),
   612 => (x"49",x"6e",x"87",x"d4"),
   613 => (x"c1",x"81",x"c8",x"c1"),
   614 => (x"c8",x"49",x"6e",x"79"),
   615 => (x"c5",x"4c",x"69",x"81"),
   616 => (x"fe",x"49",x"75",x"87"),
   617 => (x"d0",x"ff",x"87",x"d7"),
   618 => (x"78",x"e1",x"c8",x"48"),
   619 => (x"48",x"74",x"7b",x"dd"),
   620 => (x"70",x"98",x"ff",x"c3"),
   621 => (x"c8",x"49",x"74",x"7b"),
   622 => (x"48",x"71",x"29",x"b7"),
   623 => (x"70",x"98",x"ff",x"c3"),
   624 => (x"d0",x"49",x"74",x"7b"),
   625 => (x"48",x"71",x"29",x"b7"),
   626 => (x"70",x"98",x"ff",x"c3"),
   627 => (x"d8",x"48",x"74",x"7b"),
   628 => (x"7b",x"70",x"28",x"b7"),
   629 => (x"7b",x"7b",x"7b",x"c0"),
   630 => (x"7b",x"7b",x"7b",x"7b"),
   631 => (x"7b",x"7b",x"7b",x"7b"),
   632 => (x"48",x"d0",x"ff",x"7b"),
   633 => (x"75",x"78",x"e0",x"c0"),
   634 => (x"ff",x"49",x"dc",x"1e"),
   635 => (x"c4",x"87",x"e6",x"d6"),
   636 => (x"26",x"8e",x"fc",x"86"),
   637 => (x"26",x"4c",x"26",x"4d"),
   638 => (x"14",x"4f",x"26",x"4b"),
   639 => (x"14",x"00",x"00",x"1d"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

