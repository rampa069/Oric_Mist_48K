library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity TEST108J is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of TEST108J is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4F",X"72",X"69",X"63",X"20",X"44",X"69",X"61",X"67",X"20",X"52",X"4F",X"4D",X"20",X"56",X"31",
		X"2E",X"30",X"38",X"6A",X"20",X"28",X"43",X"29",X"20",X"32",X"30",X"30",X"38",X"20",X"4D",X"69",
		X"6B",X"65",X"20",X"42",X"72",X"6F",X"77",X"EE",X"E6",X"02",X"40",X"48",X"AD",X"0D",X"03",X"10",
		X"07",X"8D",X"0D",X"03",X"25",X"03",X"D0",X"15",X"48",X"A2",X"00",X"A0",X"1B",X"A9",X"03",X"20",
		X"4D",X"C1",X"68",X"A0",X"1B",X"A2",X"18",X"20",X"D0",X"C4",X"4C",X"0C",X"FF",X"E6",X"00",X"D0",
		X"02",X"E6",X"01",X"68",X"40",X"78",X"D8",X"A2",X"FF",X"9A",X"A9",X"AA",X"85",X"00",X"C5",X"00",
		X"D0",X"0B",X"85",X"01",X"C5",X"01",X"D0",X"05",X"2A",X"B0",X"F1",X"90",X"03",X"4C",X"04",X"FF",
		X"E8",X"86",X"00",X"86",X"01",X"A0",X"02",X"A9",X"AA",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"08",X"FF",X"2A",X"B0",X"F4",X"C8",X"D0",X"EF",X"E6",X"01",X"A5",X"01",X"C9",X"03",X"D0",X"04",
		X"E6",X"01",X"D0",X"E3",X"C9",X"C0",X"D0",X"DF",X"20",X"9A",X"C6",X"20",X"8F",X"C5",X"20",X"A5",
		X"C5",X"20",X"1B",X"C6",X"20",X"0A",X"C1",X"20",X"2F",X"C6",X"20",X"0A",X"C1",X"20",X"9A",X"C5",
		X"20",X"BE",X"C5",X"20",X"43",X"C6",X"20",X"25",X"C6",X"20",X"0A",X"C1",X"20",X"8F",X"C5",X"20",
		X"A5",X"C5",X"20",X"61",X"C6",X"20",X"0A",X"C1",X"20",X"6B",X"C6",X"20",X"F9",X"C6",X"20",X"32",
		X"C7",X"20",X"87",X"C7",X"20",X"E0",X"C7",X"20",X"26",X"C8",X"20",X"97",X"C8",X"20",X"F4",X"C8",
		X"20",X"57",X"C6",X"20",X"0A",X"C1",X"20",X"A5",X"C5",X"20",X"42",X"CA",X"20",X"76",X"CA",X"20",
		X"40",X"CB",X"20",X"76",X"C9",X"20",X"0A",X"C1",X"20",X"AD",X"CB",X"20",X"6C",X"C9",X"20",X"0A",
		X"C1",X"20",X"A5",X"C5",X"20",X"24",X"C5",X"4C",X"00",X"FF",X"A9",X"04",X"A2",X"07",X"A0",X"1B",
		X"20",X"4D",X"C1",X"A9",X"00",X"85",X"02",X"A5",X"02",X"F0",X"FC",X"A9",X"05",X"A2",X"07",X"A0",
		X"1B",X"20",X"4D",X"C1",X"A2",X"00",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"F8",X"86",X"02",
		X"60",X"A2",X"00",X"A0",X"00",X"C4",X"08",X"D0",X"04",X"E4",X"09",X"F0",X"0F",X"B1",X"04",X"91",
		X"06",X"C8",X"D0",X"F1",X"E6",X"05",X"E6",X"07",X"E8",X"4C",X"35",X"C1",X"60",X"0A",X"69",X"93",
		X"85",X"06",X"A9",X"00",X"69",X"C1",X"85",X"07",X"98",X"48",X"A0",X"00",X"B1",X"06",X"85",X"04",
		X"C8",X"B1",X"06",X"85",X"05",X"8A",X"18",X"69",X"80",X"85",X"06",X"A9",X"00",X"69",X"BB",X"85",
		X"07",X"68",X"0A",X"0A",X"0A",X"AA",X"A0",X"05",X"18",X"65",X"06",X"85",X"06",X"90",X"02",X"E6",
		X"07",X"8A",X"88",X"D0",X"F3",X"B1",X"04",X"30",X"05",X"91",X"06",X"C8",X"D0",X"F7",X"29",X"7F",
		X"91",X"06",X"60",X"10",X"00",X"00",X"C0",X"D7",X"C1",X"EB",X"C1",X"0D",X"C2",X"27",X"C2",X"41",
		X"C2",X"8D",X"C2",X"B2",X"C2",X"D7",X"C2",X"FC",X"C2",X"05",X"C3",X"0E",X"C3",X"17",X"C3",X"24",
		X"C3",X"31",X"C3",X"3E",X"C3",X"4A",X"C3",X"5B",X"C3",X"63",X"C3",X"6F",X"C3",X"95",X"C3",X"BB",
		X"C3",X"C8",X"C3",X"D4",X"C3",X"E0",X"C3",X"EC",X"C3",X"F5",X"C3",X"1B",X"C4",X"41",X"C4",X"52",
		X"C4",X"5D",X"C4",X"68",X"C4",X"8E",X"C4",X"12",X"00",X"52",X"41",X"4D",X"20",X"54",X"65",X"73",
		X"74",X"20",X"50",X"61",X"73",X"73",X"65",X"64",X"20",X"20",X"90",X"11",X"07",X"0C",X"55",X"6E",
		X"65",X"78",X"70",X"65",X"63",X"74",X"65",X"64",X"20",X"49",X"6E",X"74",X"65",X"72",X"72",X"75",
		X"70",X"74",X"20",X"2D",X"2D",X"20",X"48",X"61",X"6C",X"74",X"65",X"64",X"A1",X"12",X"00",X"50",
		X"72",X"65",X"73",X"73",X"20",X"4E",X"4D",X"49",X"20",X"74",X"6F",X"20",X"63",X"6F",X"6E",X"74",
		X"69",X"6E",X"75",X"65",X"20",X"20",X"90",X"10",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"90",X"17",X"00",X"09",X"20",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",
		X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",
		X"3B",X"3C",X"3D",X"3E",X"3F",X"20",X"20",X"20",X"20",X"17",X"00",X"09",X"20",X"40",X"41",X"42",
		X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",
		X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"DF",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"A0",X"11",X"00",X"52",X"65",X"6D",X"6F",X"76",X"65",X"20",X"50",X"72",X"69",X"6E",X"74",
		X"65",X"72",X"20",X"4C",X"6F",X"6F",X"70",X"62",X"61",X"63",X"6B",X"20",X"43",X"6F",X"6E",X"6E",
		X"65",X"63",X"74",X"6F",X"72",X"20",X"90",X"11",X"00",X"46",X"69",X"74",X"20",X"50",X"72",X"69",
		X"6E",X"74",X"65",X"72",X"20",X"41",X"6E",X"64",X"20",X"43",X"61",X"73",X"73",X"65",X"74",X"74",
		X"65",X"20",X"4C",X"6F",X"6F",X"70",X"62",X"61",X"63",X"6B",X"20",X"90",X"12",X"00",X"50",X"41",
		X"53",X"53",X"20",X"20",X"A0",X"11",X"00",X"46",X"41",X"49",X"4C",X"20",X"20",X"A0",X"13",X"00",
		X"54",X"65",X"73",X"74",X"69",X"6E",X"E7",X"17",X"00",X"56",X"49",X"41",X"20",X"50",X"72",X"65",
		X"73",X"65",X"6E",X"F4",X"17",X"00",X"56",X"49",X"41",X"20",X"54",X"69",X"6D",X"65",X"72",X"20",
		X"B1",X"17",X"00",X"56",X"49",X"41",X"20",X"54",X"69",X"6D",X"65",X"72",X"20",X"B2",X"17",X"00",
		X"56",X"49",X"41",X"20",X"50",X"4F",X"52",X"54",X"20",X"C1",X"17",X"00",X"43",X"61",X"73",X"73",
		X"20",X"4F",X"2F",X"52",X"6C",X"79",X"2F",X"53",X"70",X"6B",X"F2",X"17",X"00",X"43",X"61",X"73",
		X"73",X"20",X"C9",X"17",X"00",X"53",X"74",X"72",X"6F",X"62",X"65",X"2F",X"41",X"63",X"EB",X"11",
		X"00",X"52",X"65",X"6D",X"6F",X"76",X"65",X"20",X"4B",X"65",X"79",X"62",X"6F",X"61",X"72",X"64",
		X"20",X"4C",X"6F",X"6F",X"70",X"62",X"61",X"63",X"6B",X"20",X"43",X"6F",X"6E",X"6E",X"65",X"63",
		X"74",X"6F",X"72",X"20",X"90",X"11",X"00",X"20",X"20",X"46",X"69",X"74",X"20",X"4B",X"65",X"79",
		X"62",X"6F",X"61",X"72",X"64",X"20",X"4C",X"6F",X"6F",X"70",X"62",X"61",X"63",X"6B",X"20",X"43",
		X"6F",X"6E",X"6E",X"65",X"63",X"74",X"6F",X"72",X"20",X"20",X"90",X"17",X"00",X"50",X"53",X"47",
		X"20",X"50",X"72",X"65",X"73",X"65",X"6E",X"F4",X"17",X"00",X"50",X"53",X"47",X"20",X"43",X"68",
		X"61",X"6E",X"20",X"C1",X"17",X"00",X"50",X"53",X"47",X"20",X"43",X"68",X"61",X"6E",X"20",X"C2",
		X"17",X"00",X"50",X"53",X"47",X"20",X"43",X"68",X"61",X"6E",X"20",X"C3",X"13",X"00",X"43",X"4F",
		X"4E",X"46",X"49",X"52",X"CD",X"13",X"00",X"43",X"6F",X"6E",X"66",X"69",X"72",X"6D",X"20",X"33",
		X"20",X"74",X"6F",X"6E",X"65",X"2F",X"6E",X"6F",X"69",X"73",X"65",X"20",X"28",X"4C",X"6F",X"20",
		X"4D",X"69",X"64",X"20",X"48",X"69",X"67",X"68",X"29",X"20",X"90",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"A0",X"17",X"00",X"50",X"53",X"47",X"20",X"50",X"6F",X"72",X"74",X"20",X"41",X"20",X"4C",X"6F",
		X"6F",X"F0",X"17",X"00",X"50",X"53",X"47",X"20",X"4E",X"6F",X"69",X"73",X"E5",X"17",X"00",X"50",
		X"53",X"47",X"20",X"53",X"77",X"65",X"65",X"F0",X"13",X"00",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"43",X"6F",X"6E",X"66",X"69",X"72",X"6D",X"20",X"74",X"6F",X"6E",X"65",X"20",
		X"73",X"77",X"65",X"65",X"70",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"90",X"12",X"00",
		X"20",X"20",X"20",X"41",X"6C",X"6C",X"20",X"74",X"65",X"73",X"74",X"73",X"20",X"70",X"61",X"73",
		X"73",X"65",X"64",X"2C",X"20",X"66",X"69",X"74",X"20",X"6B",X"65",X"79",X"62",X"6F",X"61",X"72",
		X"64",X"20",X"20",X"A0",X"85",X"0A",X"98",X"48",X"A9",X"80",X"A0",X"07",X"66",X"0A",X"69",X"30",
		X"99",X"10",X"00",X"A9",X"00",X"88",X"10",X"F4",X"68",X"A8",X"A9",X"00",X"20",X"4D",X"C1",X"60",
		X"48",X"29",X"0F",X"09",X"B0",X"C9",X"BA",X"90",X"02",X"69",X"06",X"85",X"11",X"68",X"4A",X"4A",
		X"4A",X"4A",X"09",X"30",X"C9",X"3A",X"90",X"02",X"69",X"06",X"85",X"10",X"A9",X"00",X"20",X"4D",
		X"C1",X"60",X"48",X"8A",X"48",X"98",X"48",X"BA",X"E8",X"E8",X"E8",X"BD",X"00",X"01",X"A2",X"00",
		X"A0",X"19",X"20",X"D0",X"C4",X"BA",X"E8",X"E8",X"BD",X"00",X"01",X"A2",X"03",X"A0",X"19",X"20",
		X"D0",X"C4",X"BA",X"E8",X"BD",X"00",X"01",X"A2",X"06",X"A0",X"19",X"20",X"D0",X"C4",X"68",X"A8",
		X"68",X"AA",X"68",X"60",X"A9",X"21",X"A2",X"00",X"A0",X"05",X"20",X"4D",X"C1",X"60",X"A2",X"00",
		X"A0",X"00",X"F0",X"1B",X"A5",X"0A",X"81",X"06",X"E6",X"06",X"D0",X"02",X"E6",X"07",X"A5",X"09",
		X"05",X"08",X"F0",X"0B",X"A5",X"08",X"D0",X"02",X"C6",X"09",X"C6",X"08",X"4C",X"34",X"C5",X"B1",
		X"04",X"C8",X"D0",X"02",X"E6",X"05",X"C9",X"1B",X"D0",X"15",X"B1",X"04",X"85",X"08",X"C8",X"D0",
		X"02",X"E6",X"05",X"B1",X"04",X"85",X"09",X"C8",X"D0",X"02",X"E6",X"05",X"4C",X"3E",X"C5",X"C9",
		X"19",X"D0",X"0E",X"B1",X"04",X"85",X"08",X"C8",X"D0",X"02",X"E6",X"05",X"86",X"09",X"4C",X"3E",
		X"C5",X"C9",X"1F",X"F0",X"09",X"85",X"0A",X"86",X"08",X"86",X"09",X"4C",X"34",X"C5",X"60",X"A2",
		X"05",X"20",X"E1",X"C5",X"A2",X"0B",X"20",X"E1",X"C5",X"60",X"A2",X"11",X"20",X"E1",X"C5",X"A2",
		X"17",X"20",X"E1",X"C5",X"60",X"A9",X"1A",X"8D",X"DF",X"BF",X"A9",X"20",X"8D",X"80",X"BB",X"A2",
		X"1D",X"20",X"E1",X"C5",X"A9",X"01",X"A2",X"00",X"A0",X"00",X"20",X"4D",X"C1",X"60",X"A9",X"1E",
		X"8D",X"DF",X"BF",X"A9",X"40",X"8D",X"00",X"A0",X"A2",X"23",X"20",X"E1",X"C5",X"A9",X"20",X"8D",
		X"68",X"BF",X"A2",X"29",X"20",X"E1",X"C5",X"A9",X"01",X"A2",X"01",X"A0",X"19",X"20",X"4D",X"C1",
		X"60",X"A0",X"06",X"BD",X"F1",X"C5",X"99",X"03",X"00",X"CA",X"88",X"D0",X"F6",X"20",X"31",X"C1",
		X"60",X"F5",X"CB",X"00",X"B5",X"00",X"03",X"F5",X"CE",X"00",X"B9",X"00",X"02",X"F5",X"CB",X"00",
		X"99",X"00",X"03",X"F5",X"CE",X"00",X"9D",X"00",X"02",X"80",X"BB",X"81",X"BB",X"5E",X"04",X"00",
		X"A0",X"01",X"A0",X"3F",X"1F",X"68",X"BF",X"69",X"BF",X"76",X"00",X"A9",X"02",X"A2",X"0A",X"A0",
		X"03",X"20",X"4D",X"C1",X"60",X"A9",X"06",X"A2",X"00",X"A0",X"19",X"20",X"4D",X"C1",X"60",X"A9",
		X"F5",X"85",X"04",X"A9",X"D0",X"85",X"05",X"A9",X"A8",X"85",X"06",X"A9",X"BB",X"85",X"07",X"20",
		X"2E",X"C5",X"60",X"A9",X"3A",X"85",X"04",X"A9",X"D3",X"85",X"05",X"A9",X"00",X"85",X"06",X"A9",
		X"A0",X"85",X"07",X"20",X"2E",X"C5",X"60",X"A9",X"08",X"A2",X"02",X"A0",X"02",X"20",X"4D",X"C1",
		X"60",X"A9",X"09",X"A2",X"02",X"A0",X"02",X"20",X"4D",X"C1",X"60",X"A9",X"07",X"A2",X"02",X"A0",
		X"02",X"20",X"4D",X"C1",X"60",X"A2",X"00",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"F8",X"38",
		X"E9",X"01",X"D0",X"F1",X"60",X"98",X"48",X"8A",X"48",X"A5",X"01",X"20",X"D0",X"C4",X"68",X"AA",
		X"E8",X"E8",X"68",X"A8",X"A5",X"00",X"20",X"D0",X"C4",X"60",X"A9",X"40",X"8D",X"02",X"03",X"A9",
		X"00",X"8D",X"03",X"03",X"8D",X"0B",X"03",X"8D",X"00",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A5",
		X"7F",X"8D",X"0E",X"03",X"A9",X"01",X"20",X"75",X"C6",X"A5",X"FF",X"8D",X"0D",X"03",X"60",X"09",
		X"80",X"8D",X"0E",X"03",X"29",X"7F",X"85",X"03",X"98",X"48",X"8A",X"48",X"A9",X"00",X"85",X"00",
		X"85",X"01",X"58",X"A9",X"09",X"20",X"75",X"C6",X"78",X"68",X"AA",X"68",X"A8",X"20",X"85",X"C6",
		X"60",X"A9",X"0B",X"A2",X"12",X"20",X"4D",X"C1",X"20",X"9A",X"C6",X"4C",X"10",X"FF",X"A9",X"0A",
		X"A2",X"12",X"20",X"4D",X"C1",X"20",X"9A",X"C6",X"60",X"A9",X"0D",X"A2",X"00",X"A0",X"04",X"20",
		X"4D",X"C1",X"A9",X"0C",X"A2",X"12",X"A0",X"04",X"20",X"4D",X"C1",X"A9",X"0F",X"8D",X"03",X"03",
		X"A2",X"0F",X"8E",X"01",X"03",X"8A",X"4D",X"01",X"03",X"29",X"0F",X"D0",X"10",X"8A",X"4D",X"0F",
		X"03",X"29",X"0F",X"D0",X"08",X"CA",X"10",X"EA",X"A0",X"04",X"4C",X"EE",X"C6",X"A0",X"04",X"4C",
		X"E1",X"C6",X"A9",X"0E",X"A2",X"00",X"A0",X"05",X"20",X"4D",X"C1",X"A9",X"0C",X"A2",X"12",X"A0",
		X"05",X"20",X"4D",X"C1",X"A9",X"40",X"8D",X"0B",X"03",X"A9",X"10",X"8D",X"04",X"03",X"A9",X"27",
		X"8D",X"05",X"03",X"A9",X"40",X"A0",X"05",X"A2",X"1E",X"20",X"C6",X"C6",X"A5",X"00",X"D0",X"22",
		X"A5",X"01",X"D0",X"1E",X"A9",X"40",X"A0",X"05",X"A2",X"23",X"20",X"BF",X"C6",X"A5",X"01",X"C9",
		X"01",X"D0",X"0F",X"A5",X"00",X"C9",X"26",X"30",X"09",X"C9",X"2E",X"10",X"05",X"A0",X"05",X"4C",
		X"EE",X"C6",X"A0",X"05",X"4C",X"E1",X"C6",X"A9",X"0F",X"A2",X"00",X"A0",X"06",X"20",X"4D",X"C1",
		X"A9",X"0C",X"A2",X"12",X"A0",X"06",X"20",X"4D",X"C1",X"A9",X"00",X"8D",X"0B",X"03",X"A9",X"00",
		X"8D",X"08",X"03",X"A9",X"FA",X"8D",X"09",X"03",X"A9",X"20",X"A0",X"06",X"A2",X"1E",X"20",X"C6",
		X"C6",X"A5",X"00",X"D0",X"26",X"A5",X"01",X"D0",X"22",X"A9",X"00",X"8D",X"08",X"03",X"A9",X"FA",
		X"8D",X"09",X"03",X"A9",X"20",X"A0",X"06",X"A2",X"23",X"20",X"BF",X"C6",X"A5",X"01",X"D0",X"0B",
		X"A5",X"00",X"C9",X"01",X"D0",X"05",X"A0",X"06",X"4C",X"EE",X"C6",X"A0",X"06",X"4C",X"E1",X"C6",
		X"A9",X"10",X"A2",X"00",X"A0",X"07",X"20",X"4D",X"C1",X"A9",X"F0",X"8D",X"03",X"03",X"A2",X"0F",
		X"8A",X"0A",X"0A",X"0A",X"0A",X"8D",X"01",X"03",X"8A",X"4D",X"01",X"03",X"29",X"0F",X"D0",X"21",
		X"CA",X"10",X"ED",X"A9",X"0F",X"8D",X"03",X"03",X"A2",X"0F",X"8E",X"01",X"03",X"8A",X"0A",X"0A",
		X"0A",X"0A",X"4D",X"01",X"03",X"29",X"F0",X"D0",X"08",X"CA",X"10",X"EE",X"A0",X"07",X"4C",X"EE",
		X"C6",X"A0",X"07",X"4C",X"E1",X"C6",X"A9",X"11",X"A2",X"00",X"A0",X"08",X"20",X"4D",X"C1",X"A9",
		X"0C",X"A2",X"12",X"A0",X"08",X"20",X"4D",X"C1",X"A9",X"04",X"A2",X"07",X"A0",X"1B",X"20",X"4D",
		X"C1",X"A9",X"C0",X"8D",X"0B",X"03",X"A9",X"71",X"8D",X"04",X"03",X"A9",X"02",X"8D",X"05",X"03",
		X"A9",X"40",X"8D",X"02",X"03",X"A9",X"14",X"85",X"0B",X"A9",X"40",X"8D",X"00",X"03",X"A9",X"01",
		X"20",X"75",X"C6",X"A5",X"02",X"D0",X"14",X"A9",X"00",X"8D",X"00",X"03",X"A9",X"01",X"20",X"75",
		X"C6",X"A5",X"02",X"D0",X"06",X"C6",X"0B",X"D0",X"E0",X"F0",X"0E",X"A9",X"05",X"A2",X"07",X"A0",
		X"1B",X"20",X"4D",X"C1",X"A0",X"08",X"4C",X"EE",X"C6",X"A9",X"05",X"A2",X"07",X"A0",X"1B",X"20",
		X"4D",X"C1",X"A0",X"08",X"4C",X"E1",X"C6",X"A9",X"12",X"A2",X"00",X"A0",X"09",X"20",X"4D",X"C1",
		X"A9",X"0C",X"A2",X"12",X"A0",X"09",X"20",X"4D",X"C1",X"A9",X"C0",X"8D",X"0B",X"03",X"A9",X"71",
		X"8D",X"04",X"03",X"A9",X"02",X"8D",X"05",X"03",X"A9",X"40",X"8D",X"02",X"03",X"8D",X"00",X"03",
		X"A9",X"10",X"A2",X"1E",X"A0",X"09",X"20",X"C6",X"C6",X"A5",X"00",X"D0",X"22",X"A5",X"01",X"D0",
		X"1E",X"A9",X"10",X"A2",X"23",X"A0",X"09",X"20",X"BF",X"C6",X"A5",X"01",X"C9",X"09",X"D0",X"0F",
		X"A5",X"00",X"C9",X"8A",X"30",X"09",X"C9",X"99",X"10",X"05",X"A0",X"09",X"4C",X"EE",X"C6",X"A0",
		X"09",X"4C",X"E1",X"C6",X"A9",X"13",X"A2",X"00",X"A0",X"0A",X"20",X"4D",X"C1",X"A9",X"0C",X"A2",
		X"12",X"A0",X"0A",X"20",X"4D",X"C1",X"A9",X"10",X"8D",X"02",X"03",X"A9",X"00",X"8D",X"00",X"03",
		X"A9",X"01",X"8D",X"0C",X"03",X"A9",X"02",X"A0",X"0A",X"A2",X"1E",X"20",X"C6",X"C6",X"A5",X"00",
		X"D0",X"45",X"A5",X"01",X"D0",X"41",X"A9",X"82",X"8D",X"0E",X"03",X"58",X"A9",X"00",X"85",X"00",
		X"85",X"01",X"A9",X"10",X"8D",X"00",X"03",X"A9",X"01",X"20",X"75",X"C6",X"A9",X"00",X"8D",X"00",
		X"03",X"A9",X"01",X"20",X"75",X"C6",X"A9",X"10",X"8D",X"00",X"03",X"A9",X"01",X"20",X"75",X"C6",
		X"78",X"A2",X"23",X"A0",X"0A",X"20",X"85",X"C6",X"A5",X"01",X"D0",X"0B",X"A5",X"00",X"C9",X"02",
		X"D0",X"05",X"A0",X"0A",X"4C",X"EE",X"C6",X"A0",X"0A",X"4C",X"E1",X"C6",X"A9",X"14",X"A2",X"01",
		X"A0",X"02",X"20",X"4D",X"C1",X"60",X"A9",X"15",X"A2",X"01",X"A0",X"02",X"20",X"4D",X"C1",X"60",
		X"4C",X"6B",X"C6",X"08",X"48",X"78",X"A9",X"FF",X"8D",X"03",X"03",X"A9",X"CC",X"8D",X"0C",X"03",
		X"68",X"8D",X"0F",X"03",X"A8",X"8A",X"C0",X"07",X"D0",X"02",X"09",X"40",X"48",X"A9",X"EE",X"8D",
		X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"68",X"8D",X"0F",X"03",X"A9",X"EC",X"8D",X"0C",X"03",
		X"A9",X"CC",X"8D",X"0C",X"03",X"28",X"60",X"08",X"48",X"78",X"A9",X"FF",X"8D",X"03",X"03",X"A9",
		X"CC",X"8D",X"0C",X"03",X"68",X"8D",X"0F",X"03",X"A9",X"EE",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",
		X"0C",X"03",X"A9",X"00",X"8D",X"03",X"03",X"A9",X"CE",X"8D",X"0C",X"03",X"AE",X"0F",X"03",X"A9",
		X"CC",X"8D",X"0C",X"03",X"28",X"60",X"A9",X"0B",X"A2",X"12",X"20",X"4D",X"C1",X"A2",X"18",X"A0",
		X"CA",X"20",X"FF",X"C9",X"4C",X"14",X"FF",X"A9",X"0A",X"A2",X"12",X"20",X"4D",X"C1",X"60",X"08",
		X"78",X"86",X"0E",X"84",X"0F",X"A0",X"00",X"B1",X"0E",X"AA",X"98",X"48",X"20",X"83",X"C9",X"68",
		X"A8",X"C8",X"C0",X"0E",X"D0",X"F1",X"28",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"5E",X"00",X"27",X"00",X"0F",X"3F",X"0F",X"0F",
		X"0F",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"FE",X"07",X"00",X"00",X"00",
		X"00",X"00",X"A9",X"16",X"A2",X"00",X"A0",X"04",X"20",X"4D",X"C1",X"A9",X"0C",X"A2",X"12",X"A0",
		X"04",X"20",X"4D",X"C1",X"A2",X"00",X"8A",X"48",X"A9",X"00",X"20",X"83",X"C9",X"A9",X"00",X"20",
		X"B7",X"C9",X"68",X"86",X"0A",X"45",X"0A",X"D0",X"08",X"CA",X"D0",X"EA",X"A0",X"04",X"4C",X"F7",
		X"C9",X"A0",X"04",X"4C",X"E6",X"C9",X"A2",X"26",X"A0",X"CA",X"20",X"FF",X"C9",X"A9",X"40",X"8D",
		X"02",X"03",X"A9",X"00",X"8D",X"00",X"03",X"A9",X"17",X"A2",X"00",X"A0",X"05",X"20",X"4D",X"C1",
		X"A9",X"0C",X"A2",X"12",X"A0",X"05",X"20",X"4D",X"C1",X"A9",X"07",X"A2",X"3E",X"20",X"83",X"C9",
		X"A9",X"03",X"20",X"75",X"C6",X"A0",X"05",X"A2",X"12",X"A9",X"1A",X"20",X"4D",X"C1",X"A9",X"18",
		X"A2",X"00",X"A0",X"06",X"20",X"4D",X"C1",X"A9",X"0C",X"A2",X"12",X"A0",X"06",X"20",X"4D",X"C1",
		X"A9",X"07",X"A2",X"3D",X"20",X"83",X"C9",X"A9",X"03",X"20",X"75",X"C6",X"A0",X"06",X"A2",X"12",
		X"A9",X"1A",X"20",X"4D",X"C1",X"A9",X"19",X"A2",X"00",X"A0",X"07",X"20",X"4D",X"C1",X"A9",X"0C",
		X"A2",X"12",X"A0",X"07",X"20",X"4D",X"C1",X"A9",X"07",X"A2",X"3B",X"20",X"83",X"C9",X"A9",X"03",
		X"20",X"75",X"C6",X"A0",X"07",X"A2",X"12",X"A9",X"1A",X"20",X"4D",X"C1",X"A9",X"1E",X"A2",X"00",
		X"A0",X"08",X"20",X"4D",X"C1",X"A9",X"0C",X"A2",X"12",X"A0",X"08",X"20",X"4D",X"C1",X"A9",X"07",
		X"A2",X"37",X"20",X"83",X"C9",X"A9",X"03",X"20",X"75",X"C6",X"A0",X"08",X"A2",X"12",X"A9",X"1A",
		X"20",X"4D",X"C1",X"A2",X"18",X"A0",X"CA",X"20",X"FF",X"C9",X"A9",X"1B",X"A2",X"02",X"A0",X"09",
		X"20",X"4D",X"C1",X"20",X"0A",X"C1",X"A9",X"1C",X"A2",X"02",X"A0",X"09",X"20",X"4D",X"C1",X"60",
		X"A2",X"34",X"A0",X"CA",X"20",X"FF",X"C9",X"A9",X"1F",X"A2",X"00",X"A0",X"09",X"20",X"4D",X"C1",
		X"A9",X"0C",X"A2",X"12",X"A0",X"09",X"20",X"4D",X"C1",X"A9",X"FF",X"85",X"0C",X"A9",X"08",X"85",
		X"0D",X"A9",X"00",X"A6",X"0C",X"20",X"83",X"C9",X"A9",X"01",X"A6",X"0D",X"20",X"83",X"C9",X"A2",
		X"0F",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"F8",X"A5",X"0C",X"D0",X"02",X"C6",X"0D",X"C6",
		X"0C",X"D0",X"DE",X"A5",X"0D",X"D0",X"DA",X"A2",X"18",X"A0",X"CA",X"20",X"FF",X"C9",X"A0",X"09",
		X"A2",X"12",X"A9",X"1A",X"20",X"4D",X"C1",X"A9",X"20",X"A2",X"02",X"A0",X"0A",X"20",X"4D",X"C1",
		X"20",X"0A",X"C1",X"A9",X"1C",X"A2",X"02",X"A0",X"0A",X"20",X"4D",X"C1",X"60",X"A9",X"1D",X"A2",
		X"00",X"A0",X"0A",X"20",X"4D",X"C1",X"A9",X"0C",X"A2",X"12",X"A0",X"0A",X"20",X"4D",X"C1",X"A9",
		X"00",X"8D",X"02",X"03",X"A9",X"07",X"A2",X"FF",X"20",X"83",X"C9",X"A2",X"0F",X"8A",X"48",X"0A",
		X"0A",X"0A",X"0A",X"AA",X"A9",X"0E",X"20",X"83",X"C9",X"68",X"AA",X"AD",X"00",X"03",X"29",X"0F",
		X"49",X"08",X"85",X"0A",X"E4",X"0A",X"D0",X"08",X"CA",X"10",X"E2",X"A0",X"0A",X"4C",X"F7",X"C9",
		X"A0",X"0A",X"4C",X"E6",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"08",X"08",X"00",X"08",X"00",X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"3E",
		X"14",X"3E",X"14",X"14",X"00",X"08",X"1E",X"28",X"1C",X"0A",X"3C",X"08",X"00",X"30",X"32",X"04",
		X"08",X"10",X"26",X"06",X"00",X"10",X"28",X"28",X"10",X"2A",X"24",X"1A",X"00",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"20",X"20",X"10",X"08",X"00",X"08",X"04",X"02",
		X"02",X"02",X"04",X"08",X"00",X"08",X"2A",X"1C",X"08",X"1C",X"2A",X"08",X"00",X"00",X"08",X"08",
		X"3E",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"10",X"00",X"00",X"00",
		X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"02",X"04",
		X"08",X"10",X"20",X"00",X"00",X"1C",X"22",X"26",X"2A",X"32",X"22",X"1C",X"00",X"08",X"18",X"08",
		X"08",X"08",X"08",X"1C",X"00",X"1C",X"22",X"02",X"04",X"08",X"10",X"3E",X"00",X"3E",X"02",X"04",
		X"0C",X"02",X"22",X"1C",X"00",X"04",X"0C",X"14",X"24",X"3E",X"04",X"04",X"00",X"3E",X"20",X"3C",
		X"02",X"02",X"22",X"1C",X"00",X"0C",X"10",X"20",X"3C",X"22",X"22",X"1C",X"00",X"3E",X"02",X"04",
		X"08",X"10",X"10",X"10",X"00",X"1C",X"22",X"22",X"1C",X"22",X"22",X"1C",X"00",X"1C",X"22",X"22",
		X"1E",X"02",X"04",X"18",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"08",X"08",X"10",X"04",X"08",X"10",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"3E",
		X"00",X"3E",X"00",X"00",X"00",X"10",X"08",X"04",X"02",X"04",X"08",X"10",X"00",X"1C",X"22",X"04",
		X"08",X"08",X"00",X"08",X"00",X"1C",X"22",X"2A",X"2E",X"2C",X"20",X"1E",X"00",X"08",X"14",X"22",
		X"22",X"3E",X"22",X"22",X"00",X"3C",X"22",X"22",X"3C",X"22",X"22",X"3C",X"00",X"1C",X"22",X"20",
		X"20",X"20",X"22",X"1C",X"00",X"3C",X"22",X"22",X"22",X"22",X"22",X"3C",X"00",X"3E",X"20",X"20",
		X"3C",X"20",X"20",X"3E",X"00",X"3E",X"20",X"20",X"3C",X"20",X"20",X"20",X"00",X"1E",X"20",X"20",
		X"20",X"26",X"22",X"1E",X"00",X"22",X"22",X"22",X"3E",X"22",X"22",X"22",X"00",X"1C",X"08",X"08",
		X"08",X"08",X"08",X"1C",X"00",X"02",X"02",X"02",X"02",X"02",X"22",X"1C",X"00",X"22",X"24",X"28",
		X"30",X"28",X"24",X"22",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"3E",X"00",X"22",X"36",X"2A",
		X"2A",X"22",X"22",X"22",X"00",X"22",X"22",X"32",X"2A",X"26",X"22",X"22",X"00",X"1C",X"22",X"22",
		X"22",X"22",X"22",X"1C",X"00",X"3C",X"22",X"22",X"3C",X"20",X"20",X"20",X"00",X"1C",X"22",X"22",
		X"22",X"2A",X"24",X"1A",X"00",X"3C",X"22",X"22",X"3C",X"28",X"24",X"22",X"00",X"1C",X"22",X"20",
		X"1C",X"02",X"22",X"1C",X"00",X"3E",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"22",X"22",X"22",
		X"22",X"22",X"22",X"1C",X"00",X"22",X"22",X"22",X"22",X"22",X"14",X"08",X"00",X"22",X"22",X"22",
		X"2A",X"2A",X"36",X"22",X"00",X"22",X"22",X"14",X"08",X"14",X"22",X"22",X"00",X"22",X"22",X"14",
		X"08",X"08",X"08",X"08",X"00",X"3E",X"02",X"04",X"08",X"10",X"20",X"3E",X"00",X"1E",X"10",X"10",
		X"10",X"10",X"10",X"1E",X"00",X"00",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"3C",X"04",X"04",
		X"04",X"04",X"04",X"3C",X"00",X"08",X"14",X"2A",X"08",X"08",X"08",X"08",X"00",X"0E",X"10",X"10",
		X"10",X"3C",X"10",X"3E",X"00",X"0C",X"12",X"2D",X"29",X"29",X"2D",X"12",X"0C",X"00",X"00",X"1C",
		X"02",X"1E",X"22",X"1E",X"00",X"20",X"20",X"3C",X"22",X"22",X"22",X"3C",X"00",X"00",X"00",X"1E",
		X"20",X"20",X"20",X"1E",X"00",X"02",X"02",X"1E",X"22",X"22",X"22",X"1E",X"00",X"00",X"00",X"1C",
		X"22",X"3E",X"20",X"1E",X"00",X"0C",X"12",X"10",X"3C",X"10",X"10",X"10",X"00",X"00",X"00",X"1C",
		X"22",X"22",X"1E",X"02",X"1C",X"20",X"20",X"3C",X"22",X"22",X"22",X"22",X"00",X"08",X"00",X"18",
		X"08",X"08",X"08",X"1C",X"00",X"04",X"00",X"0C",X"04",X"04",X"04",X"24",X"18",X"20",X"20",X"22",
		X"24",X"38",X"24",X"22",X"00",X"18",X"08",X"08",X"08",X"08",X"08",X"1C",X"00",X"00",X"00",X"36",
		X"2A",X"2A",X"2A",X"22",X"00",X"00",X"00",X"3C",X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"1C",
		X"22",X"22",X"22",X"1C",X"00",X"00",X"00",X"3C",X"22",X"22",X"3C",X"20",X"20",X"00",X"00",X"1E",
		X"22",X"22",X"1E",X"02",X"02",X"00",X"00",X"2E",X"30",X"20",X"20",X"20",X"00",X"00",X"00",X"1E",
		X"20",X"1C",X"02",X"3C",X"00",X"10",X"10",X"3C",X"10",X"10",X"12",X"0C",X"00",X"00",X"00",X"22",
		X"22",X"22",X"26",X"1A",X"00",X"00",X"00",X"22",X"22",X"22",X"14",X"08",X"00",X"00",X"00",X"22",
		X"22",X"2A",X"2A",X"36",X"00",X"00",X"00",X"22",X"14",X"08",X"14",X"22",X"00",X"00",X"00",X"22",
		X"22",X"22",X"1E",X"02",X"1C",X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"0E",X"18",X"18",
		X"30",X"18",X"18",X"0E",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"38",X"0C",X"0C",
		X"06",X"0C",X"0C",X"38",X"00",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"38",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"00",X"00",X"00",X"38",X"38",X"38",
		X"38",X"38",X"00",X"00",X"00",X"07",X"07",X"07",X"38",X"38",X"00",X"00",X"00",X"3F",X"3F",X"3F",
		X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"38",X"38",X"38",
		X"07",X"07",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"3F",X"3F",X"3F",
		X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"38",X"38",X"38",
		X"3F",X"3F",X"00",X"00",X"00",X"07",X"07",X"07",X"3F",X"3F",X"00",X"00",X"00",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"38",X"38",X"38",X"38",
		X"00",X"00",X"38",X"38",X"38",X"07",X"07",X"07",X"00",X"00",X"38",X"38",X"38",X"3F",X"3F",X"3F",
		X"00",X"00",X"38",X"38",X"38",X"00",X"00",X"00",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"38",X"38",X"38",X"38",X"38",X"07",X"07",X"07",X"38",X"38",X"38",X"38",X"38",X"3F",X"3F",X"3F",
		X"38",X"38",X"38",X"38",X"38",X"00",X"00",X"00",X"07",X"07",X"38",X"38",X"38",X"38",X"38",X"38",
		X"07",X"07",X"38",X"38",X"38",X"07",X"07",X"07",X"07",X"07",X"38",X"38",X"38",X"3F",X"3F",X"3F",
		X"07",X"07",X"38",X"38",X"38",X"00",X"00",X"00",X"3F",X"3F",X"38",X"38",X"38",X"38",X"38",X"38",
		X"3F",X"3F",X"38",X"38",X"38",X"07",X"07",X"07",X"3F",X"3F",X"38",X"38",X"38",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"38",X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"38",X"38",X"38",
		X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"07",X"07",X"07",X"3F",X"3F",X"3F",
		X"00",X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"38",X"38",X"07",X"07",X"07",X"38",X"38",X"38",
		X"38",X"38",X"07",X"07",X"07",X"07",X"07",X"07",X"38",X"38",X"07",X"07",X"07",X"3F",X"3F",X"3F",
		X"38",X"38",X"07",X"07",X"07",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"38",X"38",X"38",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"3F",X"3F",X"3F",
		X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"3F",X"3F",X"07",X"07",X"07",X"38",X"38",X"38",
		X"3F",X"3F",X"07",X"07",X"07",X"07",X"07",X"07",X"3F",X"3F",X"07",X"07",X"07",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"38",X"38",X"38",
		X"00",X"00",X"3F",X"3F",X"3F",X"07",X"07",X"07",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"38",X"38",X"3F",X"3F",X"3F",X"38",X"38",X"38",
		X"38",X"38",X"3F",X"3F",X"3F",X"07",X"07",X"07",X"38",X"38",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"38",X"38",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"07",X"07",X"3F",X"3F",X"3F",X"38",X"38",X"38",
		X"07",X"07",X"3F",X"3F",X"3F",X"07",X"07",X"07",X"07",X"07",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"07",X"07",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"38",X"38",X"38",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"07",X"07",X"07",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"17",X"00",X"20",X"19",X"0A",X"54",X"65",X"78",X"74",X"20",X"54",
		X"65",X"73",X"74",X"20",X"43",X"61",X"72",X"64",X"20",X"19",X"0C",X"10",X"19",X"04",X"11",X"19",
		X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",
		X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",
		X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",
		X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",
		X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",
		X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",
		X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",
		X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",
		X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",
		X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",
		X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",
		X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"05",X"00",X"20",X"19",X"25",X"17",
		X"00",X"20",X"20",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",
		X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",
		X"3D",X"3E",X"3F",X"20",X"19",X"03",X"17",X"00",X"20",X"20",X"40",X"41",X"42",X"43",X"44",X"45",
		X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",
		X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"20",X"19",X"03",X"17",X"00",X"20",
		X"20",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",
		X"7F",X"20",X"19",X"03",X"17",X"00",X"20",X"19",X"25",X"17",X"00",X"09",X"20",X"20",X"21",X"22",
		X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",
		X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"20",X"19",X"03",
		X"17",X"00",X"20",X"19",X"25",X"17",X"00",X"09",X"20",X"40",X"41",X"42",X"43",X"44",X"45",X"46",
		X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",
		X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"20",X"19",X"03",X"17",X"00",X"18",X"20",
		X"19",X"24",X"17",X"00",X"42",X"4C",X"4B",X"10",X"01",X"52",X"45",X"44",X"10",X"02",X"47",X"52",
		X"4E",X"10",X"03",X"59",X"45",X"4C",X"10",X"04",X"42",X"4C",X"55",X"10",X"05",X"4D",X"41",X"47",
		X"10",X"06",X"43",X"59",X"41",X"10",X"07",X"57",X"48",X"54",X"97",X"80",X"C2",X"CC",X"CB",X"90",
		X"81",X"D2",X"C5",X"C4",X"90",X"82",X"C7",X"D2",X"CE",X"90",X"83",X"D9",X"C5",X"CC",X"90",X"84",
		X"C2",X"CC",X"D5",X"90",X"85",X"CD",X"C1",X"C7",X"90",X"86",X"C3",X"D9",X"C1",X"90",X"87",X"D7",
		X"C8",X"D4",X"17",X"00",X"20",X"19",X"25",X"17",X"00",X"20",X"19",X"06",X"0A",X"44",X"42",X"4C",
		X"20",X"48",X"47",X"54",X"0E",X"46",X"4C",X"41",X"53",X"48",X"0B",X"57",X"53",X"53",X"5B",X"0F",
		X"57",X"53",X"53",X"5B",X"20",X"19",X"06",X"17",X"00",X"20",X"19",X"06",X"0A",X"44",X"42",X"4C",
		X"20",X"48",X"47",X"54",X"0E",X"46",X"4C",X"41",X"53",X"48",X"0B",X"57",X"53",X"53",X"5B",X"0F",
		X"57",X"53",X"53",X"5B",X"20",X"19",X"06",X"17",X"00",X"1F",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",
		X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",
		X"19",X"04",X"10",X"19",X"04",X"11",X"19",X"04",X"12",X"19",X"04",X"13",X"19",X"04",X"14",X"19",
		X"04",X"15",X"19",X"04",X"16",X"19",X"04",X"17",X"19",X"04",X"40",X"1B",X"8F",X"01",X"17",X"00",
		X"7C",X"60",X"62",X"10",X"01",X"7C",X"7E",X"7C",X"40",X"02",X"5E",X"7C",X"62",X"40",X"03",X"62",
		X"7E",X"60",X"40",X"04",X"7C",X"60",X"62",X"40",X"05",X"62",X"48",X"5E",X"40",X"06",X"5C",X"62",
		X"48",X"40",X"07",X"62",X"62",X"7E",X"17",X"00",X"62",X"60",X"64",X"10",X"01",X"62",X"60",X"62",
		X"40",X"02",X"60",X"62",X"62",X"40",X"03",X"62",X"60",X"60",X"40",X"04",X"62",X"60",X"62",X"40",
		X"05",X"76",X"54",X"60",X"40",X"06",X"62",X"62",X"54",X"40",X"07",X"62",X"62",X"48",X"17",X"00",
		X"62",X"60",X"68",X"10",X"01",X"62",X"60",X"62",X"40",X"02",X"60",X"62",X"72",X"40",X"03",X"54",
		X"60",X"60",X"40",X"04",X"62",X"60",X"62",X"40",X"05",X"6A",X"62",X"60",X"40",X"06",X"60",X"54",
		X"62",X"40",X"07",X"62",X"62",X"48",X"17",X"00",X"7C",X"60",X"70",X"10",X"01",X"7C",X"7C",X"62",
		X"40",X"02",X"60",X"7C",X"6A",X"40",X"03",X"48",X"7C",X"60",X"40",X"04",X"7C",X"60",X"62",X"40",
		X"05",X"6A",X"62",X"60",X"40",X"06",X"60",X"48",X"62",X"40",X"07",X"6A",X"7E",X"48",X"17",X"00",
		X"62",X"60",X"68",X"10",X"01",X"68",X"60",X"62",X"40",X"02",X"66",X"68",X"66",X"40",X"03",X"48",
		X"60",X"60",X"40",X"04",X"62",X"60",X"62",X"40",X"05",X"62",X"7E",X"66",X"40",X"06",X"60",X"48",
		X"7E",X"40",X"07",X"6A",X"62",X"48",X"17",X"00",X"62",X"60",X"64",X"10",X"01",X"64",X"60",X"62",
		X"40",X"02",X"62",X"64",X"62",X"40",X"03",X"48",X"60",X"60",X"40",X"04",X"62",X"60",X"62",X"40",
		X"05",X"62",X"62",X"62",X"40",X"06",X"62",X"48",X"62",X"40",X"07",X"76",X"62",X"48",X"17",X"00",
		X"7C",X"7E",X"62",X"10",X"01",X"62",X"7E",X"7C",X"40",X"02",X"5E",X"62",X"62",X"40",X"03",X"48",
		X"7E",X"7E",X"40",X"04",X"7C",X"7E",X"5C",X"40",X"05",X"62",X"62",X"5E",X"40",X"06",X"5C",X"48",
		X"62",X"40",X"07",X"62",X"62",X"48",X"17",X"00",X"40",X"40",X"40",X"10",X"01",X"40",X"19",X"03",
		X"02",X"40",X"19",X"03",X"03",X"40",X"19",X"03",X"04",X"40",X"19",X"03",X"05",X"40",X"19",X"03",
		X"06",X"40",X"19",X"03",X"07",X"40",X"19",X"52",X"97",X"80",X"FC",X"E0",X"E2",X"90",X"81",X"FC",
		X"FE",X"FC",X"C0",X"82",X"DE",X"FC",X"E2",X"C0",X"83",X"E2",X"FE",X"E0",X"C0",X"84",X"FC",X"E0",
		X"E2",X"C0",X"85",X"E2",X"C8",X"DE",X"C0",X"86",X"DC",X"E2",X"C8",X"C0",X"87",X"E2",X"E2",X"FE",
		X"97",X"80",X"E2",X"E0",X"E4",X"90",X"81",X"E2",X"E0",X"E2",X"C0",X"82",X"E0",X"E2",X"E2",X"C0",
		X"83",X"E2",X"E0",X"E0",X"C0",X"84",X"E2",X"E0",X"E2",X"C0",X"85",X"F6",X"D4",X"E0",X"C0",X"86",
		X"E2",X"E2",X"D4",X"C0",X"87",X"E2",X"E2",X"C8",X"97",X"80",X"E2",X"E0",X"E8",X"90",X"81",X"E2",
		X"E0",X"E2",X"C0",X"82",X"E0",X"E2",X"F2",X"C0",X"83",X"D4",X"E0",X"E0",X"C0",X"84",X"E2",X"E0",
		X"E2",X"C0",X"85",X"EA",X"E2",X"E0",X"C0",X"86",X"E0",X"D4",X"E2",X"C0",X"87",X"E2",X"E2",X"C8",
		X"97",X"80",X"FC",X"E0",X"F0",X"90",X"81",X"FC",X"FC",X"E2",X"C0",X"82",X"E0",X"FC",X"EA",X"C0",
		X"83",X"C8",X"FC",X"E0",X"C0",X"84",X"FC",X"E0",X"E2",X"C0",X"85",X"EA",X"E2",X"E0",X"C0",X"86",
		X"E0",X"C8",X"E2",X"C0",X"87",X"EA",X"FE",X"C8",X"97",X"80",X"E2",X"E0",X"E8",X"90",X"81",X"E8",
		X"E0",X"E2",X"C0",X"82",X"E6",X"E8",X"E6",X"C0",X"83",X"C8",X"E0",X"E0",X"C0",X"84",X"E2",X"E0",
		X"E2",X"C0",X"85",X"E2",X"FE",X"E6",X"C0",X"86",X"E0",X"C8",X"FE",X"C0",X"87",X"EA",X"E2",X"C8",
		X"97",X"80",X"E2",X"E0",X"E4",X"90",X"81",X"E4",X"E0",X"E2",X"C0",X"82",X"E2",X"E4",X"E2",X"C0",
		X"83",X"C8",X"E0",X"E0",X"C0",X"84",X"E2",X"E0",X"E2",X"C0",X"85",X"E2",X"E2",X"E2",X"C0",X"86",
		X"E2",X"C8",X"E2",X"C0",X"87",X"F6",X"E2",X"C8",X"97",X"80",X"FC",X"FE",X"E2",X"90",X"81",X"E2",
		X"FE",X"FC",X"C0",X"82",X"DE",X"E2",X"E2",X"C0",X"83",X"C8",X"FE",X"FE",X"C0",X"84",X"FC",X"FE",
		X"DC",X"C0",X"85",X"E2",X"E2",X"DE",X"C0",X"86",X"DC",X"C8",X"E2",X"C0",X"87",X"E2",X"E2",X"C8",
		X"97",X"80",X"C0",X"C0",X"C0",X"90",X"81",X"C0",X"C0",X"C0",X"C0",X"82",X"C0",X"C0",X"C0",X"C0",
		X"83",X"C0",X"C0",X"C0",X"C0",X"84",X"C0",X"C0",X"C0",X"C0",X"85",X"C0",X"C0",X"C0",X"C0",X"86",
		X"C0",X"C0",X"C0",X"C0",X"87",X"C0",X"C0",X"C0",X"10",X"07",X"0C",X"40",X"19",X"0D",X"43",X"7A",
		X"40",X"61",X"72",X"48",X"40",X"19",X"10",X"10",X"07",X"0C",X"40",X"19",X"0D",X"42",X"42",X"41",
		X"52",X"4A",X"48",X"40",X"19",X"10",X"10",X"07",X"0C",X"40",X"19",X"0D",X"42",X"42",X"42",X"4A",
		X"42",X"48",X"40",X"19",X"10",X"10",X"07",X"0C",X"40",X"19",X"0D",X"43",X"72",X"42",X"49",X"73",
		X"78",X"40",X"19",X"10",X"10",X"07",X"0C",X"40",X"19",X"0D",X"42",X"42",X"43",X"78",X"4A",X"48",
		X"40",X"19",X"10",X"10",X"07",X"0C",X"40",X"19",X"0D",X"42",X"42",X"42",X"4A",X"4A",X"48",X"40",
		X"19",X"10",X"10",X"07",X"0C",X"40",X"19",X"0D",X"42",X"43",X"7A",X"49",X"72",X"48",X"40",X"19",
		X"10",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4C",X"00",X"FF",X"FF",X"4C",X"04",X"FF",X"FF",X"4C",X"08",X"FF",X"FF",X"4C",X"0C",X"FF",X"FF",
		X"4C",X"10",X"FF",X"FF",X"4C",X"14",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"28",X"C0",X"55",X"C0",X"2B",X"C0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
