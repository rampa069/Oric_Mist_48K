library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test109 is
 port (
   addr : in  std_logic_vector(13 downto 0);
   clk  : in  std_logic;
   data : out std_logic_vector(7 downto 0)
   );
end entity;

architecture prom of test109 is
  type rom is array(0 to 16383) of std_logic_vector(7 downto 0);
  signal rom_data: rom := (
     X"4f", X"72", X"69", X"63", X"20", X"44", X"69", X"61",
     X"67", X"20", X"52", X"4f", X"4d", X"20", X"56", X"31",
     X"2e", X"30", X"39", X"46", X"28", X"43", X"29", X"20",
     X"32", X"30", X"30", X"38", X"20", X"4d", X"69", X"6b",
     X"65", X"20", X"42", X"72", X"6f", X"77", X"ee", X"e6",
     X"02", X"40", X"48", X"ad", X"0d", X"03", X"10", X"07",
     X"8d", X"0d", X"03", X"25", X"03", X"d0", X"15", X"48",
     X"a2", X"00", X"a0", X"1b", X"a9", X"03", X"20", X"2b",
     X"c1", X"68", X"a0", X"1b", X"a2", X"18", X"20", X"ae",
     X"c4", X"4c", X"0c", X"ff", X"e6", X"00", X"d0", X"02",
     X"e6", X"01", X"68", X"40", X"78", X"d8", X"a2", X"ff",
     X"9a", X"a9", X"aa", X"85", X"00", X"c5", X"00", X"d0",
     X"0b", X"85", X"01", X"c5", X"01", X"d0", X"05", X"2a",
     X"b0", X"f1", X"90", X"03", X"4c", X"04", X"ff", X"e8",
     X"86", X"00", X"86", X"01", X"a0", X"02", X"a9", X"aa",
     X"91", X"00", X"d1", X"00", X"f0", X"03", X"4c", X"08",
     X"ff", X"2a", X"b0", X"f4", X"c8", X"d0", X"ef", X"e6",
     X"01", X"a5", X"01", X"c9", X"03", X"d0", X"04", X"e6",
     X"01", X"d0", X"e3", X"c9", X"c0", X"d0", X"df", X"20",
     X"78", X"c6", X"20", X"6d", X"c5", X"20", X"83", X"c5",
     X"20", X"f9", X"c5", X"20", X"e8", X"c0", X"20", X"0d",
     X"c6", X"20", X"e8", X"c0", X"20", X"78", X"c5", X"20",
     X"9c", X"c5", X"20", X"21", X"c6", X"20", X"03", X"c6",
     X"20", X"e8", X"c0", X"20", X"6d", X"c5", X"20", X"83",
     X"c5", X"20", X"e8", X"c0", X"20", X"d5", X"c6", X"20",
     X"0e", X"c7", X"20", X"63", X"c7", X"20", X"e8", X"c0",
     X"20", X"83", X"c5", X"20", X"1e", X"ca", X"20", X"52",
     X"ca", X"20", X"1c", X"cb", X"20", X"e8", X"c0", X"20",
     X"83", X"c5", X"20", X"02", X"c5", X"4c", X"00", X"ff",
     X"a9", X"04", X"a2", X"07", X"a0", X"1b", X"20", X"2b",
     X"c1", X"a9", X"00", X"85", X"02", X"a5", X"02", X"f0",
     X"fc", X"a9", X"05", X"a2", X"07", X"a0", X"1b", X"20",
     X"2b", X"c1", X"a2", X"00", X"a0", X"00", X"88", X"d0",
     X"fd", X"ca", X"d0", X"f8", X"86", X"02", X"60", X"a2",
     X"00", X"a0", X"00", X"c4", X"08", X"d0", X"04", X"e4",
     X"09", X"f0", X"0f", X"b1", X"04", X"91", X"06", X"c8",
     X"d0", X"f1", X"e6", X"05", X"e6", X"07", X"e8", X"4c",
     X"13", X"c1", X"60", X"0a", X"69", X"71", X"85", X"06",
     X"a9", X"00", X"69", X"c1", X"85", X"07", X"98", X"48",
     X"a0", X"00", X"b1", X"06", X"85", X"04", X"c8", X"b1",
     X"06", X"85", X"05", X"8a", X"18", X"69", X"80", X"85",
     X"06", X"a9", X"00", X"69", X"bb", X"85", X"07", X"68",
     X"0a", X"0a", X"0a", X"aa", X"a0", X"05", X"18", X"65",
     X"06", X"85", X"06", X"90", X"02", X"e6", X"07", X"8a",
     X"88", X"d0", X"f3", X"b1", X"04", X"30", X"05", X"91",
     X"06", X"c8", X"d0", X"f7", X"29", X"7f", X"91", X"06",
     X"60", X"10", X"00", X"00", X"c0", X"b5", X"c1", X"c9",
     X"c1", X"eb", X"c1", X"05", X"c2", X"1f", X"c2", X"6b",
     X"c2", X"90", X"c2", X"b5", X"c2", X"da", X"c2", X"e3",
     X"c2", X"ec", X"c2", X"f5", X"c2", X"02", X"c3", X"0f",
     X"c3", X"1c", X"c3", X"28", X"c3", X"39", X"c3", X"41",
     X"c3", X"4d", X"c3", X"73", X"c3", X"99", X"c3", X"a6",
     X"c3", X"b2", X"c3", X"be", X"c3", X"ca", X"c3", X"d3",
     X"c3", X"f9", X"c3", X"1f", X"c4", X"30", X"c4", X"3b",
     X"c4", X"46", X"c4", X"6c", X"c4", X"12", X"00", X"52",
     X"41", X"4d", X"20", X"54", X"65", X"73", X"74", X"20",
     X"50", X"61", X"73", X"73", X"65", X"64", X"20", X"20",
     X"90", X"11", X"07", X"0c", X"55", X"6e", X"65", X"78",
     X"70", X"65", X"63", X"74", X"65", X"64", X"20", X"49",
     X"6e", X"74", X"65", X"72", X"72", X"75", X"70", X"74",
     X"20", X"2d", X"2d", X"20", X"48", X"61", X"6c", X"74",
     X"65", X"64", X"a1", X"12", X"00", X"50", X"72", X"65",
     X"73", X"73", X"20", X"4e", X"4d", X"49", X"20", X"74",
     X"6f", X"20", X"63", X"6f", X"6e", X"74", X"69", X"6e",
     X"75", X"65", X"20", X"20", X"90", X"10", X"00", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"90", X"17",
     X"00", X"09", X"20", X"20", X"21", X"22", X"23", X"24",
     X"25", X"26", X"27", X"28", X"29", X"2a", X"2b", X"2c",
     X"2d", X"2e", X"2f", X"30", X"31", X"32", X"33", X"34",
     X"35", X"36", X"37", X"38", X"39", X"3a", X"3b", X"3c",
     X"3d", X"3e", X"3f", X"20", X"20", X"20", X"20", X"17",
     X"00", X"09", X"20", X"40", X"41", X"42", X"43", X"44",
     X"45", X"46", X"47", X"48", X"49", X"4a", X"4b", X"4c",
     X"4d", X"4e", X"4f", X"50", X"51", X"52", X"53", X"54",
     X"55", X"56", X"57", X"58", X"59", X"5a", X"5b", X"5c",
     X"5d", X"5e", X"df", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"a0",
     X"11", X"00", X"52", X"65", X"6d", X"6f", X"76", X"65",
     X"20", X"50", X"72", X"69", X"6e", X"74", X"65", X"72",
     X"20", X"4c", X"6f", X"6f", X"70", X"62", X"61", X"63",
     X"6b", X"20", X"43", X"6f", X"6e", X"6e", X"65", X"63",
     X"74", X"6f", X"72", X"20", X"90", X"11", X"00", X"46",
     X"69", X"74", X"20", X"50", X"72", X"69", X"6e", X"74",
     X"65", X"72", X"20", X"41", X"6e", X"64", X"20", X"43",
     X"61", X"73", X"73", X"65", X"74", X"74", X"65", X"20",
     X"4c", X"6f", X"6f", X"70", X"62", X"61", X"63", X"6b",
     X"20", X"90", X"12", X"00", X"50", X"41", X"53", X"53",
     X"20", X"20", X"a0", X"11", X"00", X"46", X"41", X"49",
     X"4c", X"20", X"20", X"a0", X"13", X"00", X"54", X"65",
     X"73", X"74", X"69", X"6e", X"e7", X"17", X"00", X"56",
     X"49", X"41", X"20", X"50", X"72", X"65", X"73", X"65",
     X"6e", X"f4", X"17", X"00", X"56", X"49", X"41", X"20",
     X"54", X"69", X"6d", X"65", X"72", X"20", X"b1", X"17",
     X"00", X"56", X"49", X"41", X"20", X"54", X"69", X"6d",
     X"65", X"72", X"20", X"b2", X"17", X"00", X"56", X"49",
     X"41", X"20", X"50", X"4f", X"52", X"54", X"20", X"c1",
     X"17", X"00", X"43", X"61", X"73", X"73", X"20", X"4f",
     X"2f", X"52", X"6c", X"79", X"2f", X"53", X"70", X"6b",
     X"f2", X"17", X"00", X"43", X"61", X"73", X"73", X"20",
     X"c9", X"17", X"00", X"53", X"74", X"72", X"6f", X"62",
     X"65", X"2f", X"41", X"63", X"eb", X"11", X"00", X"52",
     X"65", X"6d", X"6f", X"76", X"65", X"20", X"4b", X"65",
     X"79", X"62", X"6f", X"61", X"72", X"64", X"20", X"4c",
     X"6f", X"6f", X"70", X"62", X"61", X"63", X"6b", X"20",
     X"43", X"6f", X"6e", X"6e", X"65", X"63", X"74", X"6f",
     X"72", X"20", X"90", X"11", X"00", X"20", X"20", X"46",
     X"69", X"74", X"20", X"4b", X"65", X"79", X"62", X"6f",
     X"61", X"72", X"64", X"20", X"4c", X"6f", X"6f", X"70",
     X"62", X"61", X"63", X"6b", X"20", X"43", X"6f", X"6e",
     X"6e", X"65", X"63", X"74", X"6f", X"72", X"20", X"20",
     X"90", X"17", X"00", X"50", X"53", X"47", X"20", X"50",
     X"72", X"65", X"73", X"65", X"6e", X"f4", X"17", X"00",
     X"50", X"53", X"47", X"20", X"43", X"68", X"61", X"6e",
     X"20", X"c1", X"17", X"00", X"50", X"53", X"47", X"20",
     X"43", X"68", X"61", X"6e", X"20", X"c2", X"17", X"00",
     X"50", X"53", X"47", X"20", X"43", X"68", X"61", X"6e",
     X"20", X"c3", X"13", X"00", X"43", X"4f", X"4e", X"46",
     X"49", X"52", X"cd", X"13", X"00", X"43", X"6f", X"6e",
     X"66", X"69", X"72", X"6d", X"20", X"33", X"20", X"74",
     X"6f", X"6e", X"65", X"2f", X"6e", X"6f", X"69", X"73",
     X"65", X"20", X"28", X"4c", X"6f", X"20", X"4d", X"69",
     X"64", X"20", X"48", X"69", X"67", X"68", X"29", X"20",
     X"90", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"a0", X"17",
     X"00", X"50", X"53", X"47", X"20", X"50", X"6f", X"72",
     X"74", X"20", X"41", X"20", X"4c", X"6f", X"6f", X"f0",
     X"17", X"00", X"50", X"53", X"47", X"20", X"4e", X"6f",
     X"69", X"73", X"e5", X"17", X"00", X"50", X"53", X"47",
     X"20", X"53", X"77", X"65", X"65", X"f0", X"13", X"00",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"43", X"6f", X"6e", X"66", X"69", X"72", X"6d",
     X"20", X"74", X"6f", X"6e", X"65", X"20", X"73", X"77",
     X"65", X"65", X"70", X"20", X"20", X"20", X"20", X"20",
     X"20", X"20", X"20", X"90", X"12", X"00", X"20", X"20",
     X"20", X"41", X"6c", X"6c", X"20", X"74", X"65", X"73",
     X"74", X"73", X"20", X"70", X"61", X"73", X"73", X"65",
     X"64", X"2c", X"20", X"66", X"69", X"74", X"20", X"6b",
     X"65", X"79", X"62", X"6f", X"61", X"72", X"64", X"20",
     X"20", X"a0", X"85", X"0a", X"98", X"48", X"a9", X"80",
     X"a0", X"07", X"66", X"0a", X"69", X"30", X"99", X"10",
     X"00", X"a9", X"00", X"88", X"10", X"f4", X"68", X"a8",
     X"a9", X"00", X"20", X"2b", X"c1", X"60", X"48", X"29",
     X"0f", X"09", X"b0", X"c9", X"ba", X"90", X"02", X"69",
     X"06", X"85", X"11", X"68", X"4a", X"4a", X"4a", X"4a",
     X"09", X"30", X"c9", X"3a", X"90", X"02", X"69", X"06",
     X"85", X"10", X"a9", X"00", X"20", X"2b", X"c1", X"60",
     X"48", X"8a", X"48", X"98", X"48", X"ba", X"e8", X"e8",
     X"e8", X"bd", X"00", X"01", X"a2", X"00", X"a0", X"19",
     X"20", X"ae", X"c4", X"ba", X"e8", X"e8", X"bd", X"00",
     X"01", X"a2", X"03", X"a0", X"19", X"20", X"ae", X"c4",
     X"ba", X"e8", X"bd", X"00", X"01", X"a2", X"06", X"a0",
     X"19", X"20", X"ae", X"c4", X"68", X"a8", X"68", X"aa",
     X"68", X"60", X"a9", X"21", X"a2", X"00", X"a0", X"05",
     X"20", X"2b", X"c1", X"60", X"a2", X"00", X"a0", X"00",
     X"f0", X"1b", X"a5", X"0a", X"81", X"06", X"e6", X"06",
     X"d0", X"02", X"e6", X"07", X"a5", X"09", X"05", X"08",
     X"f0", X"0b", X"a5", X"08", X"d0", X"02", X"c6", X"09",
     X"c6", X"08", X"4c", X"12", X"c5", X"b1", X"04", X"c8",
     X"d0", X"02", X"e6", X"05", X"c9", X"1b", X"d0", X"15",
     X"b1", X"04", X"85", X"08", X"c8", X"d0", X"02", X"e6",
     X"05", X"b1", X"04", X"85", X"09", X"c8", X"d0", X"02",
     X"e6", X"05", X"4c", X"1c", X"c5", X"c9", X"19", X"d0",
     X"0e", X"b1", X"04", X"85", X"08", X"c8", X"d0", X"02",
     X"e6", X"05", X"86", X"09", X"4c", X"1c", X"c5", X"c9",
     X"1f", X"f0", X"09", X"85", X"0a", X"86", X"08", X"86",
     X"09", X"4c", X"12", X"c5", X"60", X"a2", X"05", X"20",
     X"bf", X"c5", X"a2", X"0b", X"20", X"bf", X"c5", X"60",
     X"a2", X"11", X"20", X"bf", X"c5", X"a2", X"17", X"20",
     X"bf", X"c5", X"60", X"a9", X"1a", X"8d", X"df", X"bf",
     X"a9", X"20", X"8d", X"80", X"bb", X"a2", X"1d", X"20",
     X"bf", X"c5", X"a9", X"01", X"a2", X"00", X"a0", X"00",
     X"20", X"2b", X"c1", X"60", X"a9", X"1e", X"8d", X"df",
     X"bf", X"a9", X"40", X"8d", X"00", X"a0", X"a2", X"23",
     X"20", X"bf", X"c5", X"a9", X"20", X"8d", X"68", X"bf",
     X"a2", X"29", X"20", X"bf", X"c5", X"a9", X"01", X"a2",
     X"01", X"a0", X"19", X"20", X"2b", X"c1", X"60", X"a0",
     X"06", X"bd", X"cf", X"c5", X"99", X"03", X"00", X"ca",
     X"88", X"d0", X"f6", X"20", X"0f", X"c1", X"60", X"d1",
     X"cb", X"00", X"b5", X"00", X"03", X"d1", X"ce", X"00",
     X"b9", X"00", X"02", X"d1", X"cb", X"00", X"99", X"00",
     X"03", X"d1", X"ce", X"00", X"9d", X"00", X"02", X"80",
     X"bb", X"81", X"bb", X"5e", X"04", X"00", X"a0", X"01",
     X"a0", X"3f", X"1f", X"68", X"bf", X"69", X"bf", X"76",
     X"00", X"a9", X"02", X"a2", X"0a", X"a0", X"03", X"20",
     X"2b", X"c1", X"60", X"a9", X"06", X"a2", X"00", X"a0",
     X"19", X"20", X"2b", X"c1", X"60", X"a9", X"d1", X"85",
     X"04", X"a9", X"d0", X"85", X"05", X"a9", X"a8", X"85",
     X"06", X"a9", X"bb", X"85", X"07", X"20", X"0c", X"c5",
     X"60", X"a9", X"16", X"85", X"04", X"a9", X"d3", X"85",
     X"05", X"a9", X"00", X"85", X"06", X"a9", X"a0", X"85",
     X"07", X"20", X"0c", X"c5", X"60", X"a9", X"08", X"a2",
     X"02", X"a0", X"02", X"20", X"2b", X"c1", X"60", X"a9",
     X"09", X"a2", X"02", X"a0", X"02", X"20", X"2b", X"c1",
     X"60", X"a9", X"07", X"a2", X"02", X"a0", X"02", X"20",
     X"2b", X"c1", X"60", X"a2", X"00", X"a0", X"00", X"88",
     X"d0", X"fd", X"ca", X"d0", X"f8", X"38", X"e9", X"01",
     X"d0", X"f1", X"60", X"98", X"48", X"8a", X"48", X"a5",
     X"01", X"20", X"ae", X"c4", X"68", X"aa", X"e8", X"e8",
     X"68", X"a8", X"a5", X"00", X"20", X"ae", X"c4", X"60",
     X"a9", X"40", X"8d", X"02", X"03", X"a9", X"00", X"8d",
     X"03", X"03", X"8d", X"0b", X"03", X"8d", X"00", X"03",
     X"a9", X"cc", X"8d", X"0c", X"03", X"a5", X"7f", X"8d",
     X"0e", X"03", X"a9", X"01", X"20", X"53", X"c6", X"a5",
     X"ff", X"8d", X"0d", X"03", X"60", X"09", X"80", X"8d",
     X"0e", X"03", X"29", X"7f", X"85", X"03", X"98", X"48",
     X"8a", X"48", X"a9", X"00", X"85", X"00", X"85", X"01",
     X"58", X"a9", X"09", X"20", X"53", X"c6", X"78", X"68",
     X"aa", X"68", X"a8", X"20", X"63", X"c6", X"60", X"a9",
     X"0b", X"a2", X"12", X"20", X"2b", X"c1", X"20", X"78",
     X"c6", X"60", X"a9", X"0a", X"a2", X"12", X"20", X"2b",
     X"c1", X"20", X"78", X"c6", X"60", X"a9", X"0d", X"a2",
     X"00", X"a0", X"04", X"20", X"2b", X"c1", X"a9", X"0c",
     X"a2", X"12", X"a0", X"04", X"20", X"2b", X"c1", X"a9",
     X"0f", X"8d", X"03", X"03", X"a2", X"0f", X"8e", X"01",
     X"03", X"8a", X"4d", X"01", X"03", X"29", X"0f", X"d0",
     X"10", X"8a", X"4d", X"0f", X"03", X"29", X"0f", X"d0",
     X"08", X"ca", X"10", X"ea", X"a0", X"04", X"4c", X"ca",
     X"c6", X"a0", X"04", X"4c", X"bf", X"c6", X"a9", X"0e",
     X"a2", X"00", X"a0", X"05", X"20", X"2b", X"c1", X"a9",
     X"0c", X"a2", X"12", X"a0", X"05", X"20", X"2b", X"c1",
     X"a9", X"40", X"8d", X"0b", X"03", X"a9", X"10", X"8d",
     X"04", X"03", X"a9", X"27", X"8d", X"05", X"03", X"a9",
     X"40", X"a0", X"05", X"a2", X"1e", X"20", X"a4", X"c6",
     X"a5", X"00", X"d0", X"22", X"a5", X"01", X"d0", X"1e",
     X"a9", X"40", X"a0", X"05", X"a2", X"23", X"20", X"9d",
     X"c6", X"a5", X"01", X"c9", X"01", X"d0", X"0f", X"a5",
     X"00", X"c9", X"26", X"30", X"09", X"c9", X"2e", X"10",
     X"05", X"a0", X"05", X"4c", X"ca", X"c6", X"a0", X"05",
     X"4c", X"bf", X"c6", X"a9", X"0f", X"a2", X"00", X"a0",
     X"06", X"20", X"2b", X"c1", X"a9", X"0c", X"a2", X"12",
     X"a0", X"06", X"20", X"2b", X"c1", X"a9", X"00", X"8d",
     X"0b", X"03", X"a9", X"00", X"8d", X"08", X"03", X"a9",
     X"fa", X"8d", X"09", X"03", X"a9", X"20", X"a0", X"06",
     X"a2", X"1e", X"20", X"a4", X"c6", X"a5", X"00", X"d0",
     X"26", X"a5", X"01", X"d0", X"22", X"a9", X"00", X"8d",
     X"08", X"03", X"a9", X"fa", X"8d", X"09", X"03", X"a9",
     X"20", X"a0", X"06", X"a2", X"23", X"20", X"9d", X"c6",
     X"a5", X"01", X"d0", X"0b", X"a5", X"00", X"c9", X"01",
     X"d0", X"05", X"a0", X"06", X"4c", X"ca", X"c6", X"a0",
     X"06", X"4c", X"bf", X"c6", X"a9", X"10", X"a2", X"00",
     X"a0", X"07", X"20", X"2b", X"c1", X"a9", X"f0", X"8d",
     X"03", X"03", X"a2", X"0f", X"8a", X"0a", X"0a", X"0a",
     X"0a", X"8d", X"01", X"03", X"8a", X"4d", X"01", X"03",
     X"29", X"0f", X"d0", X"21", X"ca", X"10", X"ed", X"a9",
     X"0f", X"8d", X"03", X"03", X"a2", X"0f", X"8e", X"01",
     X"03", X"8a", X"0a", X"0a", X"0a", X"0a", X"4d", X"01",
     X"03", X"29", X"f0", X"d0", X"08", X"ca", X"10", X"ee",
     X"a0", X"07", X"4c", X"ca", X"c6", X"a0", X"07", X"4c",
     X"bf", X"c6", X"a9", X"11", X"a2", X"00", X"a0", X"08",
     X"20", X"2b", X"c1", X"a9", X"0c", X"a2", X"12", X"a0",
     X"08", X"20", X"2b", X"c1", X"a9", X"04", X"a2", X"07",
     X"a0", X"1b", X"20", X"2b", X"c1", X"a9", X"c0", X"8d",
     X"0b", X"03", X"a9", X"71", X"8d", X"04", X"03", X"a9",
     X"02", X"8d", X"05", X"03", X"a9", X"40", X"8d", X"02",
     X"03", X"a9", X"14", X"85", X"0b", X"a9", X"40", X"8d",
     X"00", X"03", X"a9", X"01", X"20", X"53", X"c6", X"a5",
     X"02", X"d0", X"14", X"a9", X"00", X"8d", X"00", X"03",
     X"a9", X"01", X"20", X"53", X"c6", X"a5", X"02", X"d0",
     X"06", X"c6", X"0b", X"d0", X"e0", X"f0", X"0e", X"a9",
     X"05", X"a2", X"07", X"a0", X"1b", X"20", X"2b", X"c1",
     X"a0", X"08", X"4c", X"ca", X"c6", X"a9", X"05", X"a2",
     X"07", X"a0", X"1b", X"20", X"2b", X"c1", X"a0", X"08",
     X"4c", X"bf", X"c6", X"a9", X"12", X"a2", X"00", X"a0",
     X"09", X"20", X"2b", X"c1", X"a9", X"0c", X"a2", X"12",
     X"a0", X"09", X"20", X"2b", X"c1", X"a9", X"c0", X"8d",
     X"0b", X"03", X"a9", X"71", X"8d", X"04", X"03", X"a9",
     X"02", X"8d", X"05", X"03", X"a9", X"40", X"8d", X"02",
     X"03", X"8d", X"00", X"03", X"a9", X"10", X"a2", X"1e",
     X"a0", X"09", X"20", X"a4", X"c6", X"a5", X"00", X"d0",
     X"22", X"a5", X"01", X"d0", X"1e", X"a9", X"10", X"a2",
     X"23", X"a0", X"09", X"20", X"9d", X"c6", X"a5", X"01",
     X"c9", X"09", X"d0", X"0f", X"a5", X"00", X"c9", X"8a",
     X"30", X"09", X"c9", X"99", X"10", X"05", X"a0", X"09",
     X"4c", X"ca", X"c6", X"a0", X"09", X"4c", X"bf", X"c6",
     X"a9", X"13", X"a2", X"00", X"a0", X"0a", X"20", X"2b",
     X"c1", X"a9", X"0c", X"a2", X"12", X"a0", X"0a", X"20",
     X"2b", X"c1", X"a9", X"10", X"8d", X"02", X"03", X"a9",
     X"00", X"8d", X"00", X"03", X"a9", X"01", X"8d", X"0c",
     X"03", X"a9", X"02", X"a0", X"0a", X"a2", X"1e", X"20",
     X"a4", X"c6", X"a5", X"00", X"d0", X"45", X"a5", X"01",
     X"d0", X"41", X"a9", X"82", X"8d", X"0e", X"03", X"58",
     X"a9", X"00", X"85", X"00", X"85", X"01", X"a9", X"10",
     X"8d", X"00", X"03", X"a9", X"01", X"20", X"53", X"c6",
     X"a9", X"00", X"8d", X"00", X"03", X"a9", X"01", X"20",
     X"53", X"c6", X"a9", X"10", X"8d", X"00", X"03", X"a9",
     X"01", X"20", X"53", X"c6", X"78", X"a2", X"23", X"a0",
     X"0a", X"20", X"63", X"c6", X"a5", X"01", X"d0", X"0b",
     X"a5", X"00", X"c9", X"02", X"d0", X"05", X"a0", X"0a",
     X"4c", X"ca", X"c6", X"a0", X"0a", X"4c", X"bf", X"c6",
     X"a9", X"14", X"a2", X"01", X"a0", X"02", X"20", X"2b",
     X"c1", X"60", X"a9", X"15", X"a2", X"01", X"a0", X"02",
     X"20", X"2b", X"c1", X"60", X"4c", X"49", X"c6", X"08",
     X"48", X"78", X"a9", X"ff", X"8d", X"03", X"03", X"a9",
     X"cc", X"8d", X"0c", X"03", X"68", X"8d", X"0f", X"03",
     X"a8", X"8a", X"c0", X"07", X"d0", X"02", X"09", X"40",
     X"48", X"a9", X"ee", X"8d", X"0c", X"03", X"a9", X"cc",
     X"8d", X"0c", X"03", X"68", X"8d", X"0f", X"03", X"a9",
     X"ec", X"8d", X"0c", X"03", X"a9", X"cc", X"8d", X"0c",
     X"03", X"28", X"60", X"08", X"48", X"78", X"a9", X"ff",
     X"8d", X"03", X"03", X"a9", X"cc", X"8d", X"0c", X"03",
     X"68", X"8d", X"0f", X"03", X"a9", X"ee", X"8d", X"0c",
     X"03", X"a9", X"cc", X"8d", X"0c", X"03", X"a9", X"00",
     X"8d", X"03", X"03", X"a9", X"ce", X"8d", X"0c", X"03",
     X"ae", X"0f", X"03", X"a9", X"cc", X"8d", X"0c", X"03",
     X"28", X"60", X"a9", X"0b", X"a2", X"12", X"20", X"2b",
     X"c1", X"a2", X"f4", X"a0", X"c9", X"20", X"db", X"c9",
     X"4c", X"14", X"ff", X"a9", X"0a", X"a2", X"12", X"20",
     X"2b", X"c1", X"60", X"08", X"78", X"86", X"0e", X"84",
     X"0f", X"a0", X"00", X"b1", X"0e", X"aa", X"98", X"48",
     X"20", X"5f", X"c9", X"68", X"a8", X"c8", X"c0", X"0e",
     X"d0", X"f1", X"28", X"60", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"3f", X"00", X"00", X"00", X"00",
     X"00", X"00", X"ee", X"00", X"5e", X"00", X"27", X"00",
     X"0f", X"3f", X"0f", X"0f", X"0f", X"00", X"00", X"00",
     X"ff", X"0f", X"00", X"00", X"00", X"00", X"00", X"fe",
     X"07", X"00", X"00", X"00", X"00", X"00", X"a9", X"16",
     X"a2", X"00", X"a0", X"04", X"20", X"2b", X"c1", X"a9",
     X"0c", X"a2", X"12", X"a0", X"04", X"20", X"2b", X"c1",
     X"a2", X"00", X"8a", X"48", X"a9", X"00", X"20", X"5f",
     X"c9", X"a9", X"00", X"20", X"93", X"c9", X"68", X"86",
     X"0a", X"45", X"0a", X"d0", X"08", X"ca", X"d0", X"ea",
     X"a0", X"04", X"4c", X"d3", X"c9", X"a0", X"04", X"4c",
     X"c2", X"c9", X"a2", X"02", X"a0", X"ca", X"20", X"db",
     X"c9", X"a9", X"40", X"8d", X"02", X"03", X"a9", X"00",
     X"8d", X"00", X"03", X"a9", X"17", X"a2", X"00", X"a0",
     X"05", X"20", X"2b", X"c1", X"a9", X"0c", X"a2", X"12",
     X"a0", X"05", X"20", X"2b", X"c1", X"a9", X"07", X"a2",
     X"3e", X"20", X"5f", X"c9", X"a9", X"03", X"20", X"53",
     X"c6", X"a0", X"05", X"a2", X"12", X"a9", X"1a", X"20",
     X"2b", X"c1", X"a9", X"18", X"a2", X"00", X"a0", X"06",
     X"20", X"2b", X"c1", X"a9", X"0c", X"a2", X"12", X"a0",
     X"06", X"20", X"2b", X"c1", X"a9", X"07", X"a2", X"3d",
     X"20", X"5f", X"c9", X"a9", X"03", X"20", X"53", X"c6",
     X"a0", X"06", X"a2", X"12", X"a9", X"1a", X"20", X"2b",
     X"c1", X"a9", X"19", X"a2", X"00", X"a0", X"07", X"20",
     X"2b", X"c1", X"a9", X"0c", X"a2", X"12", X"a0", X"07",
     X"20", X"2b", X"c1", X"a9", X"07", X"a2", X"3b", X"20",
     X"5f", X"c9", X"a9", X"03", X"20", X"53", X"c6", X"a0",
     X"07", X"a2", X"12", X"a9", X"1a", X"20", X"2b", X"c1",
     X"a9", X"1e", X"a2", X"00", X"a0", X"08", X"20", X"2b",
     X"c1", X"a9", X"0c", X"a2", X"12", X"a0", X"08", X"20",
     X"2b", X"c1", X"a9", X"07", X"a2", X"37", X"20", X"5f",
     X"c9", X"a9", X"03", X"20", X"53", X"c6", X"a0", X"08",
     X"a2", X"12", X"a9", X"1a", X"20", X"2b", X"c1", X"a2",
     X"f4", X"a0", X"c9", X"20", X"db", X"c9", X"a9", X"1b",
     X"a2", X"02", X"a0", X"09", X"20", X"2b", X"c1", X"20",
     X"e8", X"c0", X"a9", X"1c", X"a2", X"02", X"a0", X"09",
     X"20", X"2b", X"c1", X"60", X"a2", X"10", X"a0", X"ca",
     X"20", X"db", X"c9", X"a9", X"1f", X"a2", X"00", X"a0",
     X"09", X"20", X"2b", X"c1", X"a9", X"0c", X"a2", X"12",
     X"a0", X"09", X"20", X"2b", X"c1", X"a9", X"ff", X"85",
     X"0c", X"a9", X"08", X"85", X"0d", X"a9", X"00", X"a6",
     X"0c", X"20", X"5f", X"c9", X"a9", X"01", X"a6", X"0d",
     X"20", X"5f", X"c9", X"a2", X"0f", X"a0", X"00", X"88",
     X"d0", X"fd", X"ca", X"d0", X"f8", X"a5", X"0c", X"d0",
     X"02", X"c6", X"0d", X"c6", X"0c", X"d0", X"de", X"a5",
     X"0d", X"d0", X"da", X"a2", X"f4", X"a0", X"c9", X"20",
     X"db", X"c9", X"a0", X"09", X"a2", X"12", X"a9", X"1a",
     X"20", X"2b", X"c1", X"a9", X"20", X"a2", X"02", X"a0",
     X"0a", X"20", X"2b", X"c1", X"20", X"e8", X"c0", X"a9",
     X"1c", X"a2", X"02", X"a0", X"0a", X"20", X"2b", X"c1",
     X"60", X"a9", X"1d", X"a2", X"00", X"a0", X"0a", X"20",
     X"2b", X"c1", X"a9", X"0c", X"a2", X"12", X"a0", X"0a",
     X"20", X"2b", X"c1", X"a9", X"00", X"8d", X"02", X"03",
     X"a9", X"07", X"a2", X"ff", X"20", X"5f", X"c9", X"a2",
     X"0f", X"8a", X"48", X"0a", X"0a", X"0a", X"0a", X"aa",
     X"a9", X"0e", X"20", X"5f", X"c9", X"68", X"aa", X"ad",
     X"00", X"03", X"29", X"0f", X"49", X"08", X"85", X"0a",
     X"e4", X"0a", X"d0", X"08", X"ca", X"10", X"e2", X"a0",
     X"0a", X"4c", X"d3", X"c9", X"a0", X"0a", X"4c", X"c2",
     X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"08", X"08", X"08", X"08", X"08", X"00", X"08",
     X"00", X"14", X"14", X"14", X"00", X"00", X"00", X"00",
     X"00", X"14", X"14", X"3e", X"14", X"3e", X"14", X"14",
     X"00", X"08", X"1e", X"28", X"1c", X"0a", X"3c", X"08",
     X"00", X"30", X"32", X"04", X"08", X"10", X"26", X"06",
     X"00", X"10", X"28", X"28", X"10", X"2a", X"24", X"1a",
     X"00", X"08", X"08", X"08", X"00", X"00", X"00", X"00",
     X"00", X"08", X"10", X"20", X"20", X"20", X"10", X"08",
     X"00", X"08", X"04", X"02", X"02", X"02", X"04", X"08",
     X"00", X"08", X"2a", X"1c", X"08", X"1c", X"2a", X"08",
     X"00", X"00", X"08", X"08", X"3e", X"08", X"08", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"08",
     X"10", X"00", X"00", X"00", X"3e", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"00",
     X"00", X"00", X"02", X"04", X"08", X"10", X"20", X"00",
     X"00", X"1c", X"22", X"26", X"2a", X"32", X"22", X"1c",
     X"00", X"08", X"18", X"08", X"08", X"08", X"08", X"1c",
     X"00", X"1c", X"22", X"02", X"04", X"08", X"10", X"3e",
     X"00", X"3e", X"02", X"04", X"0c", X"02", X"22", X"1c",
     X"00", X"04", X"0c", X"14", X"24", X"3e", X"04", X"04",
     X"00", X"3e", X"20", X"3c", X"02", X"02", X"22", X"1c",
     X"00", X"0c", X"10", X"20", X"3c", X"22", X"22", X"1c",
     X"00", X"3e", X"02", X"04", X"08", X"10", X"10", X"10",
     X"00", X"1c", X"22", X"22", X"1c", X"22", X"22", X"1c",
     X"00", X"1c", X"22", X"22", X"1e", X"02", X"04", X"18",
     X"00", X"00", X"00", X"08", X"00", X"00", X"08", X"00",
     X"00", X"00", X"00", X"08", X"00", X"00", X"08", X"08",
     X"10", X"04", X"08", X"10", X"20", X"10", X"08", X"04",
     X"00", X"00", X"00", X"3e", X"00", X"3e", X"00", X"00",
     X"00", X"10", X"08", X"04", X"02", X"04", X"08", X"10",
     X"00", X"1c", X"22", X"04", X"08", X"08", X"00", X"08",
     X"00", X"1c", X"22", X"2a", X"2e", X"2c", X"20", X"1e",
     X"00", X"08", X"14", X"22", X"22", X"3e", X"22", X"22",
     X"00", X"3c", X"22", X"22", X"3c", X"22", X"22", X"3c",
     X"00", X"1c", X"22", X"20", X"20", X"20", X"22", X"1c",
     X"00", X"3c", X"22", X"22", X"22", X"22", X"22", X"3c",
     X"00", X"3e", X"20", X"20", X"3c", X"20", X"20", X"3e",
     X"00", X"3e", X"20", X"20", X"3c", X"20", X"20", X"20",
     X"00", X"1e", X"20", X"20", X"20", X"26", X"22", X"1e",
     X"00", X"22", X"22", X"22", X"3e", X"22", X"22", X"22",
     X"00", X"1c", X"08", X"08", X"08", X"08", X"08", X"1c",
     X"00", X"02", X"02", X"02", X"02", X"02", X"22", X"1c",
     X"00", X"22", X"24", X"28", X"30", X"28", X"24", X"22",
     X"00", X"20", X"20", X"20", X"20", X"20", X"20", X"3e",
     X"00", X"22", X"36", X"2a", X"2a", X"22", X"22", X"22",
     X"00", X"22", X"22", X"32", X"2a", X"26", X"22", X"22",
     X"00", X"1c", X"22", X"22", X"22", X"22", X"22", X"1c",
     X"00", X"3c", X"22", X"22", X"3c", X"20", X"20", X"20",
     X"00", X"1c", X"22", X"22", X"22", X"2a", X"24", X"1a",
     X"00", X"3c", X"22", X"22", X"3c", X"28", X"24", X"22",
     X"00", X"1c", X"22", X"20", X"1c", X"02", X"22", X"1c",
     X"00", X"3e", X"08", X"08", X"08", X"08", X"08", X"08",
     X"00", X"22", X"22", X"22", X"22", X"22", X"22", X"1c",
     X"00", X"22", X"22", X"22", X"22", X"22", X"14", X"08",
     X"00", X"22", X"22", X"22", X"2a", X"2a", X"36", X"22",
     X"00", X"22", X"22", X"14", X"08", X"14", X"22", X"22",
     X"00", X"22", X"22", X"14", X"08", X"08", X"08", X"08",
     X"00", X"3e", X"02", X"04", X"08", X"10", X"20", X"3e",
     X"00", X"1e", X"10", X"10", X"10", X"10", X"10", X"1e",
     X"00", X"00", X"20", X"10", X"08", X"04", X"02", X"00",
     X"00", X"3c", X"04", X"04", X"04", X"04", X"04", X"3c",
     X"00", X"08", X"14", X"2a", X"08", X"08", X"08", X"08",
     X"00", X"0e", X"10", X"10", X"10", X"3c", X"10", X"3e",
     X"00", X"0c", X"12", X"2d", X"29", X"29", X"2d", X"12",
     X"0c", X"00", X"00", X"1c", X"02", X"1e", X"22", X"1e",
     X"00", X"20", X"20", X"3c", X"22", X"22", X"22", X"3c",
     X"00", X"00", X"00", X"1e", X"20", X"20", X"20", X"1e",
     X"00", X"02", X"02", X"1e", X"22", X"22", X"22", X"1e",
     X"00", X"00", X"00", X"1c", X"22", X"3e", X"20", X"1e",
     X"00", X"0c", X"12", X"10", X"3c", X"10", X"10", X"10",
     X"00", X"00", X"00", X"1c", X"22", X"22", X"1e", X"02",
     X"1c", X"20", X"20", X"3c", X"22", X"22", X"22", X"22",
     X"00", X"08", X"00", X"18", X"08", X"08", X"08", X"1c",
     X"00", X"04", X"00", X"0c", X"04", X"04", X"04", X"24",
     X"18", X"20", X"20", X"22", X"24", X"38", X"24", X"22",
     X"00", X"18", X"08", X"08", X"08", X"08", X"08", X"1c",
     X"00", X"00", X"00", X"36", X"2a", X"2a", X"2a", X"22",
     X"00", X"00", X"00", X"3c", X"22", X"22", X"22", X"22",
     X"00", X"00", X"00", X"1c", X"22", X"22", X"22", X"1c",
     X"00", X"00", X"00", X"3c", X"22", X"22", X"3c", X"20",
     X"20", X"00", X"00", X"1e", X"22", X"22", X"1e", X"02",
     X"02", X"00", X"00", X"2e", X"30", X"20", X"20", X"20",
     X"00", X"00", X"00", X"1e", X"20", X"1c", X"02", X"3c",
     X"00", X"10", X"10", X"3c", X"10", X"10", X"12", X"0c",
     X"00", X"00", X"00", X"22", X"22", X"22", X"26", X"1a",
     X"00", X"00", X"00", X"22", X"22", X"22", X"14", X"08",
     X"00", X"00", X"00", X"22", X"22", X"2a", X"2a", X"36",
     X"00", X"00", X"00", X"22", X"14", X"08", X"14", X"22",
     X"00", X"00", X"00", X"22", X"22", X"22", X"1e", X"02",
     X"1c", X"00", X"00", X"3e", X"04", X"08", X"10", X"3e",
     X"00", X"0e", X"18", X"18", X"30", X"18", X"18", X"0e",
     X"00", X"08", X"08", X"08", X"08", X"08", X"08", X"08",
     X"08", X"38", X"0c", X"0c", X"06", X"0c", X"0c", X"38",
     X"00", X"2a", X"15", X"2a", X"15", X"2a", X"15", X"2a",
     X"15", X"3f", X"3f", X"3f", X"3f", X"3f", X"3f", X"3f",
     X"3f", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"38", X"38", X"38", X"00", X"00", X"00", X"00",
     X"00", X"07", X"07", X"07", X"00", X"00", X"00", X"00",
     X"00", X"3f", X"3f", X"3f", X"00", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"38", X"38", X"00", X"00",
     X"00", X"38", X"38", X"38", X"38", X"38", X"00", X"00",
     X"00", X"07", X"07", X"07", X"38", X"38", X"00", X"00",
     X"00", X"3f", X"3f", X"3f", X"38", X"38", X"00", X"00",
     X"00", X"00", X"00", X"00", X"07", X"07", X"00", X"00",
     X"00", X"38", X"38", X"38", X"07", X"07", X"00", X"00",
     X"00", X"07", X"07", X"07", X"07", X"07", X"00", X"00",
     X"00", X"3f", X"3f", X"3f", X"07", X"07", X"00", X"00",
     X"00", X"00", X"00", X"00", X"3f", X"3f", X"00", X"00",
     X"00", X"38", X"38", X"38", X"3f", X"3f", X"00", X"00",
     X"00", X"07", X"07", X"07", X"3f", X"3f", X"00", X"00",
     X"00", X"3f", X"3f", X"3f", X"3f", X"3f", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"38", X"38",
     X"38", X"38", X"38", X"38", X"00", X"00", X"38", X"38",
     X"38", X"07", X"07", X"07", X"00", X"00", X"38", X"38",
     X"38", X"3f", X"3f", X"3f", X"00", X"00", X"38", X"38",
     X"38", X"00", X"00", X"00", X"38", X"38", X"38", X"38",
     X"38", X"38", X"38", X"38", X"38", X"38", X"38", X"38",
     X"38", X"07", X"07", X"07", X"38", X"38", X"38", X"38",
     X"38", X"3f", X"3f", X"3f", X"38", X"38", X"38", X"38",
     X"38", X"00", X"00", X"00", X"07", X"07", X"38", X"38",
     X"38", X"38", X"38", X"38", X"07", X"07", X"38", X"38",
     X"38", X"07", X"07", X"07", X"07", X"07", X"38", X"38",
     X"38", X"3f", X"3f", X"3f", X"07", X"07", X"38", X"38",
     X"38", X"00", X"00", X"00", X"3f", X"3f", X"38", X"38",
     X"38", X"38", X"38", X"38", X"3f", X"3f", X"38", X"38",
     X"38", X"07", X"07", X"07", X"3f", X"3f", X"38", X"38",
     X"38", X"3f", X"3f", X"3f", X"3f", X"3f", X"38", X"38",
     X"38", X"00", X"00", X"00", X"00", X"00", X"07", X"07",
     X"07", X"38", X"38", X"38", X"00", X"00", X"07", X"07",
     X"07", X"07", X"07", X"07", X"00", X"00", X"07", X"07",
     X"07", X"3f", X"3f", X"3f", X"00", X"00", X"07", X"07",
     X"07", X"00", X"00", X"00", X"38", X"38", X"07", X"07",
     X"07", X"38", X"38", X"38", X"38", X"38", X"07", X"07",
     X"07", X"07", X"07", X"07", X"38", X"38", X"07", X"07",
     X"07", X"3f", X"3f", X"3f", X"38", X"38", X"07", X"07",
     X"07", X"00", X"00", X"00", X"07", X"07", X"07", X"07",
     X"07", X"38", X"38", X"38", X"07", X"07", X"07", X"07",
     X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07",
     X"07", X"3f", X"3f", X"3f", X"07", X"07", X"07", X"07",
     X"07", X"00", X"00", X"00", X"3f", X"3f", X"07", X"07",
     X"07", X"38", X"38", X"38", X"3f", X"3f", X"07", X"07",
     X"07", X"07", X"07", X"07", X"3f", X"3f", X"07", X"07",
     X"07", X"3f", X"3f", X"3f", X"3f", X"3f", X"07", X"07",
     X"07", X"00", X"00", X"00", X"00", X"00", X"3f", X"3f",
     X"3f", X"38", X"38", X"38", X"00", X"00", X"3f", X"3f",
     X"3f", X"07", X"07", X"07", X"00", X"00", X"3f", X"3f",
     X"3f", X"3f", X"3f", X"3f", X"00", X"00", X"3f", X"3f",
     X"3f", X"00", X"00", X"00", X"38", X"38", X"3f", X"3f",
     X"3f", X"38", X"38", X"38", X"38", X"38", X"3f", X"3f",
     X"3f", X"07", X"07", X"07", X"38", X"38", X"3f", X"3f",
     X"3f", X"3f", X"3f", X"3f", X"38", X"38", X"3f", X"3f",
     X"3f", X"00", X"00", X"00", X"07", X"07", X"3f", X"3f",
     X"3f", X"38", X"38", X"38", X"07", X"07", X"3f", X"3f",
     X"3f", X"07", X"07", X"07", X"07", X"07", X"3f", X"3f",
     X"3f", X"3f", X"3f", X"3f", X"07", X"07", X"3f", X"3f",
     X"3f", X"00", X"00", X"00", X"3f", X"3f", X"3f", X"3f",
     X"3f", X"38", X"38", X"38", X"3f", X"3f", X"3f", X"3f",
     X"3f", X"07", X"07", X"07", X"3f", X"3f", X"3f", X"3f",
     X"3f", X"3f", X"3f", X"3f", X"3f", X"3f", X"3f", X"3f",
     X"3f", X"17", X"00", X"20", X"19", X"0a", X"54", X"65",
     X"78", X"74", X"20", X"54", X"65", X"73", X"74", X"20",
     X"43", X"61", X"72", X"64", X"20", X"19", X"0c", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"04", X"10",
     X"19", X"04", X"11", X"19", X"04", X"12", X"19", X"04",
     X"13", X"19", X"04", X"14", X"19", X"04", X"15", X"19",
     X"04", X"16", X"19", X"04", X"17", X"19", X"05", X"00",
     X"20", X"19", X"25", X"17", X"00", X"20", X"20", X"20",
     X"21", X"22", X"23", X"24", X"25", X"26", X"27", X"28",
     X"29", X"2a", X"2b", X"2c", X"2d", X"2e", X"2f", X"30",
     X"31", X"32", X"33", X"34", X"35", X"36", X"37", X"38",
     X"39", X"3a", X"3b", X"3c", X"3d", X"3e", X"3f", X"20",
     X"19", X"03", X"17", X"00", X"20", X"20", X"40", X"41",
     X"42", X"43", X"44", X"45", X"46", X"47", X"48", X"49",
     X"4a", X"4b", X"4c", X"4d", X"4e", X"4f", X"50", X"51",
     X"52", X"53", X"54", X"55", X"56", X"57", X"58", X"59",
     X"5a", X"5b", X"5c", X"5d", X"5e", X"5f", X"20", X"19",
     X"03", X"17", X"00", X"20", X"20", X"60", X"61", X"62",
     X"63", X"64", X"65", X"66", X"67", X"68", X"69", X"6a",
     X"6b", X"6c", X"6d", X"6e", X"6f", X"70", X"71", X"72",
     X"73", X"74", X"75", X"76", X"77", X"78", X"79", X"7a",
     X"7b", X"7c", X"7d", X"7e", X"7f", X"20", X"19", X"03",
     X"17", X"00", X"20", X"19", X"25", X"17", X"00", X"09",
     X"20", X"20", X"21", X"22", X"23", X"24", X"25", X"26",
     X"27", X"28", X"29", X"2a", X"2b", X"2c", X"2d", X"2e",
     X"2f", X"30", X"31", X"32", X"33", X"34", X"35", X"36",
     X"37", X"38", X"39", X"3a", X"3b", X"3c", X"3d", X"3e",
     X"3f", X"20", X"19", X"03", X"17", X"00", X"20", X"19",
     X"25", X"17", X"00", X"09", X"20", X"40", X"41", X"42",
     X"43", X"44", X"45", X"46", X"47", X"48", X"49", X"4a",
     X"4b", X"4c", X"4d", X"4e", X"4f", X"50", X"51", X"52",
     X"53", X"54", X"55", X"56", X"57", X"58", X"59", X"5a",
     X"5b", X"5c", X"5d", X"5e", X"5f", X"20", X"19", X"03",
     X"17", X"00", X"18", X"20", X"19", X"24", X"17", X"00",
     X"42", X"4c", X"4b", X"10", X"01", X"52", X"45", X"44",
     X"10", X"02", X"47", X"52", X"4e", X"10", X"03", X"59",
     X"45", X"4c", X"10", X"04", X"42", X"4c", X"55", X"10",
     X"05", X"4d", X"41", X"47", X"10", X"06", X"43", X"59",
     X"41", X"10", X"07", X"57", X"48", X"54", X"97", X"80",
     X"c2", X"cc", X"cb", X"90", X"81", X"d2", X"c5", X"c4",
     X"90", X"82", X"c7", X"d2", X"ce", X"90", X"83", X"d9",
     X"c5", X"cc", X"90", X"84", X"c2", X"cc", X"d5", X"90",
     X"85", X"cd", X"c1", X"c7", X"90", X"86", X"c3", X"d9",
     X"c1", X"90", X"87", X"d7", X"c8", X"d4", X"17", X"00",
     X"20", X"19", X"25", X"17", X"00", X"20", X"19", X"06",
     X"0a", X"44", X"42", X"4c", X"20", X"48", X"47", X"54",
     X"0e", X"46", X"4c", X"41", X"53", X"48", X"0b", X"57",
     X"53", X"53", X"5b", X"0f", X"57", X"53", X"53", X"5b",
     X"20", X"19", X"06", X"17", X"00", X"20", X"19", X"06",
     X"0a", X"44", X"42", X"4c", X"20", X"48", X"47", X"54",
     X"0e", X"46", X"4c", X"41", X"53", X"48", X"0b", X"57",
     X"53", X"53", X"5b", X"0f", X"57", X"53", X"53", X"5b",
     X"20", X"19", X"06", X"17", X"00", X"1f", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"10", X"19",
     X"04", X"11", X"19", X"04", X"12", X"19", X"04", X"13",
     X"19", X"04", X"14", X"19", X"04", X"15", X"19", X"04",
     X"16", X"19", X"04", X"17", X"19", X"04", X"40", X"1b",
     X"8f", X"01", X"17", X"00", X"7c", X"60", X"62", X"10",
     X"01", X"7c", X"7e", X"7c", X"40", X"02", X"5e", X"7c",
     X"62", X"40", X"03", X"62", X"7e", X"60", X"40", X"04",
     X"7c", X"60", X"62", X"40", X"05", X"62", X"48", X"5e",
     X"40", X"06", X"5c", X"62", X"48", X"40", X"07", X"62",
     X"62", X"7e", X"17", X"00", X"62", X"60", X"64", X"10",
     X"01", X"62", X"60", X"62", X"40", X"02", X"60", X"62",
     X"62", X"40", X"03", X"62", X"60", X"60", X"40", X"04",
     X"62", X"60", X"62", X"40", X"05", X"76", X"54", X"60",
     X"40", X"06", X"62", X"62", X"54", X"40", X"07", X"62",
     X"62", X"48", X"17", X"00", X"62", X"60", X"68", X"10",
     X"01", X"62", X"60", X"62", X"40", X"02", X"60", X"62",
     X"72", X"40", X"03", X"54", X"60", X"60", X"40", X"04",
     X"62", X"60", X"62", X"40", X"05", X"6a", X"62", X"60",
     X"40", X"06", X"60", X"54", X"62", X"40", X"07", X"62",
     X"62", X"48", X"17", X"00", X"7c", X"60", X"70", X"10",
     X"01", X"7c", X"7c", X"62", X"40", X"02", X"60", X"7c",
     X"6a", X"40", X"03", X"48", X"7c", X"60", X"40", X"04",
     X"7c", X"60", X"62", X"40", X"05", X"6a", X"62", X"60",
     X"40", X"06", X"60", X"48", X"62", X"40", X"07", X"6a",
     X"7e", X"48", X"17", X"00", X"62", X"60", X"68", X"10",
     X"01", X"68", X"60", X"62", X"40", X"02", X"66", X"68",
     X"66", X"40", X"03", X"48", X"60", X"60", X"40", X"04",
     X"62", X"60", X"62", X"40", X"05", X"62", X"7e", X"66",
     X"40", X"06", X"60", X"48", X"7e", X"40", X"07", X"6a",
     X"62", X"48", X"17", X"00", X"62", X"60", X"64", X"10",
     X"01", X"64", X"60", X"62", X"40", X"02", X"62", X"64",
     X"62", X"40", X"03", X"48", X"60", X"60", X"40", X"04",
     X"62", X"60", X"62", X"40", X"05", X"62", X"62", X"62",
     X"40", X"06", X"62", X"48", X"62", X"40", X"07", X"76",
     X"62", X"48", X"17", X"00", X"7c", X"7e", X"62", X"10",
     X"01", X"62", X"7e", X"7c", X"40", X"02", X"5e", X"62",
     X"62", X"40", X"03", X"48", X"7e", X"7e", X"40", X"04",
     X"7c", X"7e", X"5c", X"40", X"05", X"62", X"62", X"5e",
     X"40", X"06", X"5c", X"48", X"62", X"40", X"07", X"62",
     X"62", X"48", X"17", X"00", X"40", X"40", X"40", X"10",
     X"01", X"40", X"19", X"03", X"02", X"40", X"19", X"03",
     X"03", X"40", X"19", X"03", X"04", X"40", X"19", X"03",
     X"05", X"40", X"19", X"03", X"06", X"40", X"19", X"03",
     X"07", X"40", X"19", X"52", X"97", X"80", X"fc", X"e0",
     X"e2", X"90", X"81", X"fc", X"fe", X"fc", X"c0", X"82",
     X"de", X"fc", X"e2", X"c0", X"83", X"e2", X"fe", X"e0",
     X"c0", X"84", X"fc", X"e0", X"e2", X"c0", X"85", X"e2",
     X"c8", X"de", X"c0", X"86", X"dc", X"e2", X"c8", X"c0",
     X"87", X"e2", X"e2", X"fe", X"97", X"80", X"e2", X"e0",
     X"e4", X"90", X"81", X"e2", X"e0", X"e2", X"c0", X"82",
     X"e0", X"e2", X"e2", X"c0", X"83", X"e2", X"e0", X"e0",
     X"c0", X"84", X"e2", X"e0", X"e2", X"c0", X"85", X"f6",
     X"d4", X"e0", X"c0", X"86", X"e2", X"e2", X"d4", X"c0",
     X"87", X"e2", X"e2", X"c8", X"97", X"80", X"e2", X"e0",
     X"e8", X"90", X"81", X"e2", X"e0", X"e2", X"c0", X"82",
     X"e0", X"e2", X"f2", X"c0", X"83", X"d4", X"e0", X"e0",
     X"c0", X"84", X"e2", X"e0", X"e2", X"c0", X"85", X"ea",
     X"e2", X"e0", X"c0", X"86", X"e0", X"d4", X"e2", X"c0",
     X"87", X"e2", X"e2", X"c8", X"97", X"80", X"fc", X"e0",
     X"f0", X"90", X"81", X"fc", X"fc", X"e2", X"c0", X"82",
     X"e0", X"fc", X"ea", X"c0", X"83", X"c8", X"fc", X"e0",
     X"c0", X"84", X"fc", X"e0", X"e2", X"c0", X"85", X"ea",
     X"e2", X"e0", X"c0", X"86", X"e0", X"c8", X"e2", X"c0",
     X"87", X"ea", X"fe", X"c8", X"97", X"80", X"e2", X"e0",
     X"e8", X"90", X"81", X"e8", X"e0", X"e2", X"c0", X"82",
     X"e6", X"e8", X"e6", X"c0", X"83", X"c8", X"e0", X"e0",
     X"c0", X"84", X"e2", X"e0", X"e2", X"c0", X"85", X"e2",
     X"fe", X"e6", X"c0", X"86", X"e0", X"c8", X"fe", X"c0",
     X"87", X"ea", X"e2", X"c8", X"97", X"80", X"e2", X"e0",
     X"e4", X"90", X"81", X"e4", X"e0", X"e2", X"c0", X"82",
     X"e2", X"e4", X"e2", X"c0", X"83", X"c8", X"e0", X"e0",
     X"c0", X"84", X"e2", X"e0", X"e2", X"c0", X"85", X"e2",
     X"e2", X"e2", X"c0", X"86", X"e2", X"c8", X"e2", X"c0",
     X"87", X"f6", X"e2", X"c8", X"97", X"80", X"fc", X"fe",
     X"e2", X"90", X"81", X"e2", X"fe", X"fc", X"c0", X"82",
     X"de", X"e2", X"e2", X"c0", X"83", X"c8", X"fe", X"fe",
     X"c0", X"84", X"fc", X"fe", X"dc", X"c0", X"85", X"e2",
     X"e2", X"de", X"c0", X"86", X"dc", X"c8", X"e2", X"c0",
     X"87", X"e2", X"e2", X"c8", X"97", X"80", X"c0", X"c0",
     X"c0", X"90", X"81", X"c0", X"c0", X"c0", X"c0", X"82",
     X"c0", X"c0", X"c0", X"c0", X"83", X"c0", X"c0", X"c0",
     X"c0", X"84", X"c0", X"c0", X"c0", X"c0", X"85", X"c0",
     X"c0", X"c0", X"c0", X"86", X"c0", X"c0", X"c0", X"c0",
     X"87", X"c0", X"c0", X"c0", X"10", X"07", X"0c", X"40",
     X"19", X"0d", X"43", X"7a", X"40", X"61", X"72", X"48",
     X"40", X"19", X"10", X"10", X"07", X"0c", X"40", X"19",
     X"0d", X"42", X"42", X"41", X"52", X"4a", X"48", X"40",
     X"19", X"10", X"10", X"07", X"0c", X"40", X"19", X"0d",
     X"42", X"42", X"42", X"4a", X"42", X"48", X"40", X"19",
     X"10", X"10", X"07", X"0c", X"40", X"19", X"0d", X"43",
     X"72", X"42", X"49", X"73", X"78", X"40", X"19", X"10",
     X"10", X"07", X"0c", X"40", X"19", X"0d", X"42", X"42",
     X"43", X"78", X"4a", X"48", X"40", X"19", X"10", X"10",
     X"07", X"0c", X"40", X"19", X"0d", X"42", X"42", X"42",
     X"4a", X"4a", X"48", X"40", X"19", X"10", X"10", X"07",
     X"0c", X"40", X"19", X"0d", X"42", X"43", X"7a", X"49",
     X"72", X"48", X"40", X"19", X"10", X"1f", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"4c", X"00", X"ff", X"ff", X"4c", X"04", X"ff", X"ff",
     X"4c", X"08", X"ff", X"ff", X"4c", X"0c", X"ff", X"ff",
     X"4c", X"10", X"ff", X"ff", X"4c", X"14", X"ff", X"ff",
     X"00", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"27", X"c0", X"54", X"c0", X"2a", X"c0");

begin

process (clk)
  begin
    if rising_edge(clk) then
      data <= rom_data(TO_INTEGER(unsigned(addr)));
    end if;
  end process;

end architecture;
