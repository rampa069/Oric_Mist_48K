`define DEMISTIFY_PARALLEL_AUDIO 1
`define DEMISTIFY_HDMI 1
`define DEMISTIFY_ZXTRES 1
`define XILINX 1
`define VGA_8BIT 1
`define USE_CLOCK_50 1
`define NO_DIRECT_UPLOAD 1
`define I2S_AUDIO 1
`define USE_AUDIO_IN 1
`define DEMISTIFY 1
