
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"c0",x"c3",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"c4",x"c0",x"c3"),
    18 => (x"48",x"dc",x"e7",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"d9",x"e7",x"c2",x"87"),
    25 => (x"d5",x"e7",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"ed",x"c1",x"87",x"f7"),
    29 => (x"e7",x"c2",x"87",x"fc"),
    30 => (x"e7",x"c2",x"4d",x"d9"),
    31 => (x"ad",x"74",x"4c",x"d9"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"86",x"f0",x"0e",x"5d"),
    37 => (x"a6",x"c4",x"4c",x"c0"),
    38 => (x"c0",x"78",x"c0",x"48"),
    39 => (x"c0",x"4b",x"a6",x"e4"),
    40 => (x"48",x"49",x"66",x"e0"),
    41 => (x"e4",x"c0",x"80",x"c1"),
    42 => (x"7e",x"11",x"58",x"a6"),
    43 => (x"f1",x"c3",x"02",x"6e"),
    44 => (x"02",x"66",x"c4",x"87"),
    45 => (x"c4",x"87",x"c6",x"c3"),
    46 => (x"78",x"c0",x"48",x"a6"),
    47 => (x"f0",x"c0",x"4a",x"6e"),
    48 => (x"da",x"c2",x"02",x"8a"),
    49 => (x"8a",x"f3",x"c0",x"87"),
    50 => (x"87",x"db",x"c2",x"02"),
    51 => (x"dc",x"02",x"8a",x"c1"),
    52 => (x"02",x"8a",x"c8",x"87"),
    53 => (x"c4",x"87",x"c8",x"c2"),
    54 => (x"87",x"d1",x"02",x"8a"),
    55 => (x"c1",x"02",x"8a",x"c3"),
    56 => (x"8a",x"c2",x"87",x"eb"),
    57 => (x"c3",x"87",x"c6",x"02"),
    58 => (x"c9",x"c2",x"05",x"8a"),
    59 => (x"73",x"83",x"c4",x"87"),
    60 => (x"69",x"89",x"c4",x"49"),
    61 => (x"c1",x"02",x"6e",x"7e"),
    62 => (x"a6",x"c8",x"87",x"c8"),
    63 => (x"c4",x"78",x"c0",x"48"),
    64 => (x"cc",x"78",x"c0",x"80"),
    65 => (x"4a",x"6e",x"4d",x"66"),
    66 => (x"cf",x"2a",x"b7",x"dc"),
    67 => (x"c4",x"48",x"6e",x"9a"),
    68 => (x"72",x"7e",x"70",x"30"),
    69 => (x"87",x"c5",x"02",x"9a"),
    70 => (x"c1",x"48",x"a6",x"c8"),
    71 => (x"06",x"aa",x"c9",x"78"),
    72 => (x"f7",x"c0",x"87",x"c5"),
    73 => (x"c0",x"87",x"c3",x"82"),
    74 => (x"66",x"c8",x"82",x"f0"),
    75 => (x"72",x"87",x"c7",x"02"),
    76 => (x"87",x"fa",x"c1",x"49"),
    77 => (x"85",x"c1",x"84",x"c1"),
    78 => (x"04",x"ad",x"b7",x"c8"),
    79 => (x"c1",x"87",x"c7",x"ff"),
    80 => (x"f0",x"c0",x"87",x"ce"),
    81 => (x"87",x"e6",x"c1",x"49"),
    82 => (x"c3",x"c1",x"84",x"c1"),
    83 => (x"73",x"83",x"c4",x"87"),
    84 => (x"6a",x"8a",x"c4",x"4a"),
    85 => (x"87",x"f1",x"c1",x"49"),
    86 => (x"4c",x"a4",x"49",x"70"),
    87 => (x"c4",x"87",x"f1",x"c0"),
    88 => (x"78",x"c1",x"48",x"a6"),
    89 => (x"c4",x"87",x"e9",x"c0"),
    90 => (x"c4",x"4a",x"73",x"83"),
    91 => (x"c0",x"49",x"6a",x"8a"),
    92 => (x"84",x"c1",x"87",x"fc"),
    93 => (x"49",x"6e",x"87",x"da"),
    94 => (x"d3",x"87",x"f3",x"c0"),
    95 => (x"c0",x"48",x"6e",x"87"),
    96 => (x"c7",x"05",x"a8",x"e5"),
    97 => (x"48",x"a6",x"c4",x"87"),
    98 => (x"87",x"c4",x"78",x"c1"),
    99 => (x"87",x"de",x"49",x"6e"),
   100 => (x"49",x"66",x"e0",x"c0"),
   101 => (x"c0",x"80",x"c1",x"48"),
   102 => (x"11",x"58",x"a6",x"e4"),
   103 => (x"fc",x"05",x"6e",x"7e"),
   104 => (x"48",x"74",x"87",x"cf"),
   105 => (x"4d",x"26",x"8e",x"f0"),
   106 => (x"4b",x"26",x"4c",x"26"),
   107 => (x"fc",x"1e",x"4f",x"26"),
   108 => (x"ff",x"4a",x"71",x"86"),
   109 => (x"48",x"69",x"49",x"c0"),
   110 => (x"70",x"98",x"c0",x"c4"),
   111 => (x"02",x"98",x"48",x"7e"),
   112 => (x"79",x"72",x"87",x"f4"),
   113 => (x"26",x"8e",x"fc",x"48"),
   114 => (x"5b",x"5e",x"0e",x"4f"),
   115 => (x"4b",x"71",x"0e",x"5c"),
   116 => (x"4a",x"13",x"4c",x"c0"),
   117 => (x"87",x"cd",x"02",x"9a"),
   118 => (x"d1",x"ff",x"49",x"72"),
   119 => (x"13",x"84",x"c1",x"87"),
   120 => (x"f3",x"05",x"9a",x"4a"),
   121 => (x"26",x"48",x"74",x"87"),
   122 => (x"26",x"4b",x"26",x"4c"),
   123 => (x"1e",x"72",x"1e",x"4f"),
   124 => (x"48",x"12",x"1e",x"73"),
   125 => (x"87",x"ca",x"02",x"11"),
   126 => (x"98",x"df",x"c3",x"4b"),
   127 => (x"02",x"88",x"73",x"9b"),
   128 => (x"4b",x"26",x"87",x"f0"),
   129 => (x"4f",x"26",x"4a",x"26"),
   130 => (x"72",x"1e",x"73",x"1e"),
   131 => (x"04",x"8b",x"c1",x"1e"),
   132 => (x"48",x"12",x"87",x"ca"),
   133 => (x"87",x"c4",x"02",x"11"),
   134 => (x"87",x"f1",x"02",x"88"),
   135 => (x"4b",x"26",x"4a",x"26"),
   136 => (x"73",x"1e",x"4f",x"26"),
   137 => (x"a9",x"73",x"81",x"48"),
   138 => (x"12",x"87",x"c5",x"02"),
   139 => (x"87",x"f6",x"05",x"53"),
   140 => (x"73",x"1e",x"4f",x"26"),
   141 => (x"c8",x"4a",x"71",x"1e"),
   142 => (x"c1",x"49",x"4b",x"66"),
   143 => (x"02",x"99",x"71",x"8b"),
   144 => (x"48",x"12",x"87",x"cf"),
   145 => (x"78",x"08",x"d4",x"ff"),
   146 => (x"8b",x"c1",x"49",x"73"),
   147 => (x"f1",x"05",x"99",x"71"),
   148 => (x"26",x"4b",x"26",x"87"),
   149 => (x"5b",x"5e",x"0e",x"4f"),
   150 => (x"4a",x"71",x"0e",x"5c"),
   151 => (x"cc",x"4c",x"d4",x"ff"),
   152 => (x"c1",x"49",x"4b",x"66"),
   153 => (x"02",x"99",x"71",x"8b"),
   154 => (x"ff",x"c3",x"87",x"ce"),
   155 => (x"73",x"52",x"6c",x"7c"),
   156 => (x"71",x"8b",x"c1",x"49"),
   157 => (x"87",x"f2",x"05",x"99"),
   158 => (x"4b",x"26",x"4c",x"26"),
   159 => (x"73",x"1e",x"4f",x"26"),
   160 => (x"4b",x"d4",x"ff",x"1e"),
   161 => (x"6b",x"7b",x"ff",x"c3"),
   162 => (x"7b",x"ff",x"c3",x"4a"),
   163 => (x"32",x"c8",x"49",x"6b"),
   164 => (x"ff",x"c3",x"b1",x"72"),
   165 => (x"c8",x"4a",x"6b",x"7b"),
   166 => (x"c3",x"b2",x"71",x"31"),
   167 => (x"49",x"6b",x"7b",x"ff"),
   168 => (x"b1",x"72",x"32",x"c8"),
   169 => (x"4b",x"26",x"48",x"71"),
   170 => (x"5e",x"0e",x"4f",x"26"),
   171 => (x"0e",x"5d",x"5c",x"5b"),
   172 => (x"d4",x"ff",x"4d",x"71"),
   173 => (x"c3",x"48",x"75",x"4c"),
   174 => (x"7c",x"70",x"98",x"ff"),
   175 => (x"bf",x"dc",x"e7",x"c2"),
   176 => (x"d0",x"87",x"c8",x"05"),
   177 => (x"30",x"c9",x"48",x"66"),
   178 => (x"d0",x"58",x"a6",x"d4"),
   179 => (x"29",x"d8",x"49",x"66"),
   180 => (x"ff",x"c3",x"48",x"71"),
   181 => (x"d0",x"7c",x"70",x"98"),
   182 => (x"29",x"d0",x"49",x"66"),
   183 => (x"ff",x"c3",x"48",x"71"),
   184 => (x"d0",x"7c",x"70",x"98"),
   185 => (x"29",x"c8",x"49",x"66"),
   186 => (x"ff",x"c3",x"48",x"71"),
   187 => (x"d0",x"7c",x"70",x"98"),
   188 => (x"ff",x"c3",x"48",x"66"),
   189 => (x"75",x"7c",x"70",x"98"),
   190 => (x"71",x"29",x"d0",x"49"),
   191 => (x"98",x"ff",x"c3",x"48"),
   192 => (x"4b",x"6c",x"7c",x"70"),
   193 => (x"4a",x"ff",x"f0",x"c9"),
   194 => (x"05",x"ab",x"ff",x"c3"),
   195 => (x"71",x"49",x"87",x"cf"),
   196 => (x"c1",x"4b",x"6c",x"7c"),
   197 => (x"87",x"c5",x"02",x"8a"),
   198 => (x"f2",x"02",x"ab",x"71"),
   199 => (x"26",x"48",x"73",x"87"),
   200 => (x"26",x"4c",x"26",x"4d"),
   201 => (x"1e",x"4f",x"26",x"4b"),
   202 => (x"d4",x"ff",x"49",x"c0"),
   203 => (x"78",x"ff",x"c3",x"48"),
   204 => (x"c8",x"c3",x"81",x"c1"),
   205 => (x"f1",x"04",x"a9",x"b7"),
   206 => (x"0e",x"4f",x"26",x"87"),
   207 => (x"5d",x"5c",x"5b",x"5e"),
   208 => (x"f0",x"ff",x"c0",x"0e"),
   209 => (x"c1",x"4d",x"f7",x"c1"),
   210 => (x"c0",x"c0",x"c0",x"c0"),
   211 => (x"d6",x"ff",x"4b",x"c0"),
   212 => (x"df",x"f8",x"c4",x"87"),
   213 => (x"75",x"1e",x"c0",x"4c"),
   214 => (x"87",x"ce",x"fd",x"49"),
   215 => (x"a8",x"c1",x"86",x"c4"),
   216 => (x"87",x"e5",x"c0",x"05"),
   217 => (x"c3",x"48",x"d4",x"ff"),
   218 => (x"1e",x"73",x"78",x"ff"),
   219 => (x"c1",x"f0",x"e1",x"c0"),
   220 => (x"f5",x"fc",x"49",x"e9"),
   221 => (x"70",x"86",x"c4",x"87"),
   222 => (x"87",x"ca",x"05",x"98"),
   223 => (x"c3",x"48",x"d4",x"ff"),
   224 => (x"48",x"c1",x"78",x"ff"),
   225 => (x"de",x"fe",x"87",x"cb"),
   226 => (x"05",x"8c",x"c1",x"87"),
   227 => (x"c0",x"87",x"c6",x"ff"),
   228 => (x"26",x"4d",x"26",x"48"),
   229 => (x"26",x"4b",x"26",x"4c"),
   230 => (x"5b",x"5e",x"0e",x"4f"),
   231 => (x"ff",x"c0",x"0e",x"5c"),
   232 => (x"4c",x"c1",x"c1",x"f0"),
   233 => (x"c3",x"48",x"d4",x"ff"),
   234 => (x"dc",x"cf",x"78",x"ff"),
   235 => (x"87",x"d9",x"f8",x"49"),
   236 => (x"1e",x"c0",x"4b",x"d3"),
   237 => (x"f1",x"fb",x"49",x"74"),
   238 => (x"70",x"86",x"c4",x"87"),
   239 => (x"87",x"ca",x"05",x"98"),
   240 => (x"c3",x"48",x"d4",x"ff"),
   241 => (x"48",x"c1",x"78",x"ff"),
   242 => (x"da",x"fd",x"87",x"cb"),
   243 => (x"05",x"8b",x"c1",x"87"),
   244 => (x"c0",x"87",x"df",x"ff"),
   245 => (x"26",x"4c",x"26",x"48"),
   246 => (x"00",x"4f",x"26",x"4b"),
   247 => (x"00",x"44",x"4d",x"43"),
   248 => (x"43",x"48",x"44",x"53"),
   249 => (x"69",x"61",x"66",x"20"),
   250 => (x"00",x"0a",x"21",x"6c"),
   251 => (x"52",x"52",x"45",x"49"),
   252 => (x"00",x"00",x"00",x"00"),
   253 => (x"00",x"49",x"50",x"53"),
   254 => (x"74",x"69",x"72",x"57"),
   255 => (x"61",x"66",x"20",x"65"),
   256 => (x"64",x"65",x"6c",x"69"),
   257 => (x"5e",x"0e",x"00",x"0a"),
   258 => (x"0e",x"5d",x"5c",x"5b"),
   259 => (x"ff",x"4d",x"ff",x"c3"),
   260 => (x"d2",x"fc",x"4b",x"d4"),
   261 => (x"1e",x"ea",x"c6",x"87"),
   262 => (x"c1",x"f0",x"e1",x"c0"),
   263 => (x"c9",x"fa",x"49",x"c8"),
   264 => (x"c1",x"86",x"c4",x"87"),
   265 => (x"87",x"c8",x"02",x"a8"),
   266 => (x"c0",x"87",x"ee",x"fd"),
   267 => (x"87",x"e8",x"c1",x"48"),
   268 => (x"70",x"87",x"cb",x"f9"),
   269 => (x"ff",x"ff",x"cf",x"49"),
   270 => (x"a9",x"ea",x"c6",x"99"),
   271 => (x"fd",x"87",x"c8",x"02"),
   272 => (x"48",x"c0",x"87",x"d7"),
   273 => (x"75",x"87",x"d1",x"c1"),
   274 => (x"4c",x"f1",x"c0",x"7b"),
   275 => (x"70",x"87",x"ec",x"fb"),
   276 => (x"ec",x"c0",x"02",x"98"),
   277 => (x"c0",x"1e",x"c0",x"87"),
   278 => (x"fa",x"c1",x"f0",x"ff"),
   279 => (x"87",x"ca",x"f9",x"49"),
   280 => (x"98",x"70",x"86",x"c4"),
   281 => (x"75",x"87",x"da",x"05"),
   282 => (x"75",x"49",x"6b",x"7b"),
   283 => (x"75",x"7b",x"75",x"7b"),
   284 => (x"c1",x"7b",x"75",x"7b"),
   285 => (x"c4",x"02",x"99",x"c0"),
   286 => (x"db",x"48",x"c1",x"87"),
   287 => (x"d7",x"48",x"c0",x"87"),
   288 => (x"05",x"ac",x"c2",x"87"),
   289 => (x"e0",x"cf",x"87",x"ca"),
   290 => (x"87",x"fd",x"f4",x"49"),
   291 => (x"87",x"c8",x"48",x"c0"),
   292 => (x"fe",x"05",x"8c",x"c1"),
   293 => (x"48",x"c0",x"87",x"f6"),
   294 => (x"4c",x"26",x"4d",x"26"),
   295 => (x"4f",x"26",x"4b",x"26"),
   296 => (x"5c",x"5b",x"5e",x"0e"),
   297 => (x"d0",x"ff",x"0e",x"5d"),
   298 => (x"d0",x"e5",x"c0",x"4d"),
   299 => (x"c2",x"4c",x"c0",x"c1"),
   300 => (x"c1",x"48",x"dc",x"e7"),
   301 => (x"49",x"f4",x"cf",x"78"),
   302 => (x"c7",x"87",x"ce",x"f4"),
   303 => (x"f9",x"7d",x"c2",x"4b"),
   304 => (x"7d",x"c3",x"87",x"e5"),
   305 => (x"49",x"74",x"1e",x"c0"),
   306 => (x"c4",x"87",x"df",x"f7"),
   307 => (x"05",x"a8",x"c1",x"86"),
   308 => (x"c2",x"4b",x"87",x"c1"),
   309 => (x"87",x"cb",x"05",x"ab"),
   310 => (x"f3",x"49",x"ec",x"cf"),
   311 => (x"48",x"c0",x"87",x"eb"),
   312 => (x"c1",x"87",x"f6",x"c0"),
   313 => (x"d4",x"ff",x"05",x"8b"),
   314 => (x"87",x"da",x"fc",x"87"),
   315 => (x"58",x"e0",x"e7",x"c2"),
   316 => (x"cd",x"05",x"98",x"70"),
   317 => (x"c0",x"1e",x"c1",x"87"),
   318 => (x"d0",x"c1",x"f0",x"ff"),
   319 => (x"87",x"ea",x"f6",x"49"),
   320 => (x"d4",x"ff",x"86",x"c4"),
   321 => (x"78",x"ff",x"c3",x"48"),
   322 => (x"c2",x"87",x"ee",x"c4"),
   323 => (x"c2",x"58",x"e4",x"e7"),
   324 => (x"48",x"d4",x"ff",x"7d"),
   325 => (x"c1",x"78",x"ff",x"c3"),
   326 => (x"26",x"4d",x"26",x"48"),
   327 => (x"26",x"4b",x"26",x"4c"),
   328 => (x"5b",x"5e",x"0e",x"4f"),
   329 => (x"71",x"0e",x"5d",x"5c"),
   330 => (x"4c",x"ff",x"c3",x"4d"),
   331 => (x"74",x"4b",x"d4",x"ff"),
   332 => (x"48",x"d0",x"ff",x"7b"),
   333 => (x"74",x"78",x"c3",x"c4"),
   334 => (x"c0",x"1e",x"75",x"7b"),
   335 => (x"d8",x"c1",x"f0",x"ff"),
   336 => (x"87",x"e6",x"f5",x"49"),
   337 => (x"98",x"70",x"86",x"c4"),
   338 => (x"cf",x"87",x"cb",x"02"),
   339 => (x"f8",x"f1",x"49",x"f8"),
   340 => (x"c0",x"48",x"c1",x"87"),
   341 => (x"7b",x"74",x"87",x"ee"),
   342 => (x"c8",x"7b",x"fe",x"c3"),
   343 => (x"66",x"d4",x"1e",x"c0"),
   344 => (x"87",x"ce",x"f3",x"49"),
   345 => (x"7b",x"74",x"86",x"c4"),
   346 => (x"7b",x"74",x"7b",x"74"),
   347 => (x"4a",x"e0",x"da",x"d8"),
   348 => (x"05",x"6b",x"7b",x"74"),
   349 => (x"8a",x"c1",x"87",x"c5"),
   350 => (x"74",x"87",x"f5",x"05"),
   351 => (x"48",x"d0",x"ff",x"7b"),
   352 => (x"48",x"c0",x"78",x"c2"),
   353 => (x"4c",x"26",x"4d",x"26"),
   354 => (x"4f",x"26",x"4b",x"26"),
   355 => (x"5c",x"5b",x"5e",x"0e"),
   356 => (x"86",x"fc",x"0e",x"5d"),
   357 => (x"d4",x"ff",x"4b",x"71"),
   358 => (x"c5",x"7e",x"c0",x"4c"),
   359 => (x"4a",x"df",x"cd",x"ee"),
   360 => (x"6c",x"7c",x"ff",x"c3"),
   361 => (x"a8",x"fe",x"c3",x"48"),
   362 => (x"87",x"f8",x"c0",x"05"),
   363 => (x"9b",x"73",x"4d",x"74"),
   364 => (x"d4",x"87",x"cc",x"02"),
   365 => (x"49",x"73",x"1e",x"66"),
   366 => (x"c4",x"87",x"da",x"f2"),
   367 => (x"ff",x"87",x"d4",x"86"),
   368 => (x"d1",x"c4",x"48",x"d0"),
   369 => (x"4a",x"66",x"d4",x"78"),
   370 => (x"c1",x"7d",x"ff",x"c3"),
   371 => (x"87",x"f8",x"05",x"8a"),
   372 => (x"c3",x"5a",x"a6",x"d8"),
   373 => (x"73",x"7c",x"7c",x"ff"),
   374 => (x"87",x"c5",x"05",x"9b"),
   375 => (x"d0",x"48",x"d0",x"ff"),
   376 => (x"7e",x"4a",x"c1",x"78"),
   377 => (x"fe",x"05",x"8a",x"c1"),
   378 => (x"48",x"6e",x"87",x"f6"),
   379 => (x"4d",x"26",x"8e",x"fc"),
   380 => (x"4b",x"26",x"4c",x"26"),
   381 => (x"73",x"1e",x"4f",x"26"),
   382 => (x"c0",x"4a",x"71",x"1e"),
   383 => (x"48",x"d4",x"ff",x"4b"),
   384 => (x"ff",x"78",x"ff",x"c3"),
   385 => (x"c3",x"c4",x"48",x"d0"),
   386 => (x"48",x"d4",x"ff",x"78"),
   387 => (x"72",x"78",x"ff",x"c3"),
   388 => (x"f0",x"ff",x"c0",x"1e"),
   389 => (x"f2",x"49",x"d1",x"c1"),
   390 => (x"86",x"c4",x"87",x"d0"),
   391 => (x"d2",x"05",x"98",x"70"),
   392 => (x"1e",x"c0",x"c8",x"87"),
   393 => (x"fd",x"49",x"66",x"cc"),
   394 => (x"86",x"c4",x"87",x"e2"),
   395 => (x"d0",x"ff",x"4b",x"70"),
   396 => (x"73",x"78",x"c2",x"48"),
   397 => (x"26",x"4b",x"26",x"48"),
   398 => (x"5b",x"5e",x"0e",x"4f"),
   399 => (x"c0",x"0e",x"5d",x"5c"),
   400 => (x"f0",x"ff",x"c0",x"1e"),
   401 => (x"f1",x"49",x"c9",x"c1"),
   402 => (x"1e",x"d2",x"87",x"e0"),
   403 => (x"49",x"ec",x"e7",x"c2"),
   404 => (x"c8",x"87",x"f9",x"fc"),
   405 => (x"c1",x"4c",x"c0",x"86"),
   406 => (x"ac",x"b7",x"d2",x"84"),
   407 => (x"c2",x"87",x"f8",x"04"),
   408 => (x"bf",x"97",x"ec",x"e7"),
   409 => (x"99",x"c0",x"c3",x"49"),
   410 => (x"05",x"a9",x"c0",x"c1"),
   411 => (x"c2",x"87",x"e7",x"c0"),
   412 => (x"bf",x"97",x"f3",x"e7"),
   413 => (x"c2",x"31",x"d0",x"49"),
   414 => (x"bf",x"97",x"f4",x"e7"),
   415 => (x"72",x"32",x"c8",x"4a"),
   416 => (x"f5",x"e7",x"c2",x"b1"),
   417 => (x"b1",x"4a",x"bf",x"97"),
   418 => (x"ff",x"cf",x"4c",x"71"),
   419 => (x"c1",x"9c",x"ff",x"ff"),
   420 => (x"c1",x"34",x"ca",x"84"),
   421 => (x"e7",x"c2",x"87",x"e7"),
   422 => (x"49",x"bf",x"97",x"f5"),
   423 => (x"99",x"c6",x"31",x"c1"),
   424 => (x"97",x"f6",x"e7",x"c2"),
   425 => (x"b7",x"c7",x"4a",x"bf"),
   426 => (x"c2",x"b1",x"72",x"2a"),
   427 => (x"bf",x"97",x"f1",x"e7"),
   428 => (x"9d",x"cf",x"4d",x"4a"),
   429 => (x"97",x"f2",x"e7",x"c2"),
   430 => (x"9a",x"c3",x"4a",x"bf"),
   431 => (x"e7",x"c2",x"32",x"ca"),
   432 => (x"4b",x"bf",x"97",x"f3"),
   433 => (x"b2",x"73",x"33",x"c2"),
   434 => (x"97",x"f4",x"e7",x"c2"),
   435 => (x"c0",x"c3",x"4b",x"bf"),
   436 => (x"2b",x"b7",x"c6",x"9b"),
   437 => (x"81",x"c2",x"b2",x"73"),
   438 => (x"30",x"71",x"48",x"c1"),
   439 => (x"48",x"c1",x"49",x"70"),
   440 => (x"4d",x"70",x"30",x"75"),
   441 => (x"84",x"c1",x"4c",x"72"),
   442 => (x"c0",x"c8",x"94",x"71"),
   443 => (x"cc",x"06",x"ad",x"b7"),
   444 => (x"b7",x"34",x"c1",x"87"),
   445 => (x"b7",x"c0",x"c8",x"2d"),
   446 => (x"f4",x"ff",x"01",x"ad"),
   447 => (x"26",x"48",x"74",x"87"),
   448 => (x"26",x"4c",x"26",x"4d"),
   449 => (x"0e",x"4f",x"26",x"4b"),
   450 => (x"5d",x"5c",x"5b",x"5e"),
   451 => (x"c2",x"86",x"fc",x"0e"),
   452 => (x"c0",x"48",x"d4",x"f0"),
   453 => (x"cc",x"e8",x"c2",x"78"),
   454 => (x"fb",x"49",x"c0",x"1e"),
   455 => (x"86",x"c4",x"87",x"d8"),
   456 => (x"c5",x"05",x"98",x"70"),
   457 => (x"c9",x"48",x"c0",x"87"),
   458 => (x"4d",x"c0",x"87",x"d5"),
   459 => (x"48",x"d0",x"f5",x"c2"),
   460 => (x"e9",x"c2",x"78",x"c1"),
   461 => (x"e6",x"c0",x"4a",x"c2"),
   462 => (x"4b",x"c8",x"49",x"d8"),
   463 => (x"70",x"87",x"c9",x"eb"),
   464 => (x"87",x"c6",x"05",x"98"),
   465 => (x"48",x"d0",x"f5",x"c2"),
   466 => (x"e9",x"c2",x"78",x"c0"),
   467 => (x"e6",x"c0",x"4a",x"de"),
   468 => (x"4b",x"c8",x"49",x"e4"),
   469 => (x"70",x"87",x"f1",x"ea"),
   470 => (x"87",x"c6",x"05",x"98"),
   471 => (x"48",x"d0",x"f5",x"c2"),
   472 => (x"f5",x"c2",x"78",x"c0"),
   473 => (x"c0",x"02",x"bf",x"d0"),
   474 => (x"ef",x"c2",x"87",x"fe"),
   475 => (x"c2",x"4d",x"bf",x"d2"),
   476 => (x"bf",x"9f",x"ca",x"f0"),
   477 => (x"c5",x"48",x"6e",x"7e"),
   478 => (x"05",x"a8",x"ea",x"d6"),
   479 => (x"ef",x"c2",x"87",x"c7"),
   480 => (x"ce",x"4d",x"bf",x"d2"),
   481 => (x"ca",x"48",x"6e",x"87"),
   482 => (x"02",x"a8",x"d5",x"e9"),
   483 => (x"48",x"c0",x"87",x"c5"),
   484 => (x"c2",x"87",x"ec",x"c7"),
   485 => (x"75",x"1e",x"cc",x"e8"),
   486 => (x"87",x"da",x"f9",x"49"),
   487 => (x"98",x"70",x"86",x"c4"),
   488 => (x"c0",x"87",x"c5",x"05"),
   489 => (x"87",x"d7",x"c7",x"48"),
   490 => (x"4a",x"de",x"e9",x"c2"),
   491 => (x"49",x"f0",x"e6",x"c0"),
   492 => (x"d3",x"e9",x"4b",x"c8"),
   493 => (x"05",x"98",x"70",x"87"),
   494 => (x"c2",x"87",x"c8",x"c0"),
   495 => (x"c1",x"48",x"d4",x"f0"),
   496 => (x"c2",x"87",x"d8",x"78"),
   497 => (x"c0",x"4a",x"c2",x"e9"),
   498 => (x"c8",x"49",x"fc",x"e6"),
   499 => (x"87",x"f8",x"e8",x"4b"),
   500 => (x"c0",x"02",x"98",x"70"),
   501 => (x"48",x"c0",x"87",x"c5"),
   502 => (x"c2",x"87",x"e4",x"c6"),
   503 => (x"bf",x"97",x"ca",x"f0"),
   504 => (x"a9",x"d5",x"c1",x"49"),
   505 => (x"87",x"cd",x"c0",x"05"),
   506 => (x"97",x"cb",x"f0",x"c2"),
   507 => (x"ea",x"c2",x"49",x"bf"),
   508 => (x"c5",x"c0",x"02",x"a9"),
   509 => (x"c6",x"48",x"c0",x"87"),
   510 => (x"e8",x"c2",x"87",x"c5"),
   511 => (x"7e",x"bf",x"97",x"cc"),
   512 => (x"e9",x"c3",x"48",x"6e"),
   513 => (x"ce",x"c0",x"02",x"a8"),
   514 => (x"c3",x"48",x"6e",x"87"),
   515 => (x"c0",x"02",x"a8",x"eb"),
   516 => (x"48",x"c0",x"87",x"c5"),
   517 => (x"c2",x"87",x"e8",x"c5"),
   518 => (x"bf",x"97",x"d7",x"e8"),
   519 => (x"c0",x"05",x"99",x"49"),
   520 => (x"e8",x"c2",x"87",x"cc"),
   521 => (x"49",x"bf",x"97",x"d8"),
   522 => (x"c0",x"02",x"a9",x"c2"),
   523 => (x"48",x"c0",x"87",x"c5"),
   524 => (x"c2",x"87",x"cc",x"c5"),
   525 => (x"bf",x"97",x"d9",x"e8"),
   526 => (x"d0",x"f0",x"c2",x"48"),
   527 => (x"48",x"4c",x"70",x"58"),
   528 => (x"f0",x"c2",x"88",x"c1"),
   529 => (x"e8",x"c2",x"58",x"d4"),
   530 => (x"49",x"bf",x"97",x"da"),
   531 => (x"e8",x"c2",x"81",x"75"),
   532 => (x"4a",x"bf",x"97",x"db"),
   533 => (x"a1",x"72",x"32",x"c8"),
   534 => (x"ec",x"f4",x"c2",x"7e"),
   535 => (x"c2",x"78",x"6e",x"48"),
   536 => (x"bf",x"97",x"dc",x"e8"),
   537 => (x"c4",x"f5",x"c2",x"48"),
   538 => (x"d4",x"f0",x"c2",x"58"),
   539 => (x"d3",x"c2",x"02",x"bf"),
   540 => (x"de",x"e9",x"c2",x"87"),
   541 => (x"cc",x"e6",x"c0",x"4a"),
   542 => (x"e6",x"4b",x"c8",x"49"),
   543 => (x"98",x"70",x"87",x"ca"),
   544 => (x"87",x"c5",x"c0",x"02"),
   545 => (x"f6",x"c3",x"48",x"c0"),
   546 => (x"cc",x"f0",x"c2",x"87"),
   547 => (x"f5",x"c2",x"4c",x"bf"),
   548 => (x"e8",x"c2",x"5c",x"c0"),
   549 => (x"49",x"bf",x"97",x"f1"),
   550 => (x"e8",x"c2",x"31",x"c8"),
   551 => (x"4a",x"bf",x"97",x"f0"),
   552 => (x"e8",x"c2",x"49",x"a1"),
   553 => (x"4a",x"bf",x"97",x"f2"),
   554 => (x"a1",x"72",x"32",x"d0"),
   555 => (x"f3",x"e8",x"c2",x"49"),
   556 => (x"d8",x"4a",x"bf",x"97"),
   557 => (x"49",x"a1",x"72",x"32"),
   558 => (x"59",x"c8",x"f5",x"c2"),
   559 => (x"bf",x"c0",x"f5",x"c2"),
   560 => (x"ec",x"f4",x"c2",x"91"),
   561 => (x"f4",x"c2",x"81",x"bf"),
   562 => (x"e8",x"c2",x"59",x"f4"),
   563 => (x"4a",x"bf",x"97",x"f9"),
   564 => (x"e8",x"c2",x"32",x"c8"),
   565 => (x"4b",x"bf",x"97",x"f8"),
   566 => (x"e8",x"c2",x"4a",x"a2"),
   567 => (x"4b",x"bf",x"97",x"fa"),
   568 => (x"a2",x"73",x"33",x"d0"),
   569 => (x"fb",x"e8",x"c2",x"4a"),
   570 => (x"cf",x"4b",x"bf",x"97"),
   571 => (x"73",x"33",x"d8",x"9b"),
   572 => (x"f4",x"c2",x"4a",x"a2"),
   573 => (x"8a",x"c2",x"5a",x"f8"),
   574 => (x"f4",x"c2",x"92",x"74"),
   575 => (x"a1",x"72",x"48",x"f8"),
   576 => (x"87",x"c7",x"c1",x"78"),
   577 => (x"97",x"de",x"e8",x"c2"),
   578 => (x"31",x"c8",x"49",x"bf"),
   579 => (x"97",x"dd",x"e8",x"c2"),
   580 => (x"49",x"a1",x"4a",x"bf"),
   581 => (x"ff",x"c7",x"31",x"c5"),
   582 => (x"c2",x"29",x"c9",x"81"),
   583 => (x"c2",x"59",x"c0",x"f5"),
   584 => (x"bf",x"97",x"e3",x"e8"),
   585 => (x"c2",x"32",x"c8",x"4a"),
   586 => (x"bf",x"97",x"e2",x"e8"),
   587 => (x"c2",x"4a",x"a2",x"4b"),
   588 => (x"c2",x"5a",x"c8",x"f5"),
   589 => (x"92",x"bf",x"c0",x"f5"),
   590 => (x"f4",x"c2",x"82",x"6e"),
   591 => (x"f4",x"c2",x"5a",x"fc"),
   592 => (x"78",x"c0",x"48",x"f4"),
   593 => (x"48",x"f0",x"f4",x"c2"),
   594 => (x"c2",x"78",x"a1",x"72"),
   595 => (x"c2",x"48",x"c8",x"f5"),
   596 => (x"78",x"bf",x"f4",x"f4"),
   597 => (x"48",x"cc",x"f5",x"c2"),
   598 => (x"bf",x"f8",x"f4",x"c2"),
   599 => (x"d4",x"f0",x"c2",x"78"),
   600 => (x"c9",x"c0",x"02",x"bf"),
   601 => (x"c4",x"48",x"74",x"87"),
   602 => (x"c0",x"7e",x"70",x"30"),
   603 => (x"f4",x"c2",x"87",x"c9"),
   604 => (x"c4",x"48",x"bf",x"fc"),
   605 => (x"c2",x"7e",x"70",x"30"),
   606 => (x"6e",x"48",x"d8",x"f0"),
   607 => (x"fc",x"48",x"c1",x"78"),
   608 => (x"26",x"4d",x"26",x"8e"),
   609 => (x"26",x"4b",x"26",x"4c"),
   610 => (x"00",x"00",x"00",x"4f"),
   611 => (x"33",x"54",x"41",x"46"),
   612 => (x"20",x"20",x"20",x"32"),
   613 => (x"00",x"00",x"00",x"00"),
   614 => (x"31",x"54",x"41",x"46"),
   615 => (x"20",x"20",x"20",x"36"),
   616 => (x"00",x"00",x"00",x"00"),
   617 => (x"33",x"54",x"41",x"46"),
   618 => (x"20",x"20",x"20",x"32"),
   619 => (x"00",x"00",x"00",x"00"),
   620 => (x"33",x"54",x"41",x"46"),
   621 => (x"20",x"20",x"20",x"32"),
   622 => (x"00",x"00",x"00",x"00"),
   623 => (x"31",x"54",x"41",x"46"),
   624 => (x"20",x"20",x"20",x"36"),
   625 => (x"5b",x"5e",x"0e",x"00"),
   626 => (x"71",x"0e",x"5d",x"5c"),
   627 => (x"d4",x"f0",x"c2",x"4a"),
   628 => (x"87",x"cb",x"02",x"bf"),
   629 => (x"2b",x"c7",x"4b",x"72"),
   630 => (x"ff",x"c1",x"4d",x"72"),
   631 => (x"72",x"87",x"c9",x"9d"),
   632 => (x"72",x"2b",x"c8",x"4b"),
   633 => (x"9d",x"ff",x"c3",x"4d"),
   634 => (x"bf",x"ec",x"f4",x"c2"),
   635 => (x"d0",x"fe",x"c0",x"83"),
   636 => (x"d9",x"02",x"ab",x"bf"),
   637 => (x"d4",x"fe",x"c0",x"87"),
   638 => (x"cc",x"e8",x"c2",x"5b"),
   639 => (x"ef",x"49",x"73",x"1e"),
   640 => (x"86",x"c4",x"87",x"f4"),
   641 => (x"c5",x"05",x"98",x"70"),
   642 => (x"c0",x"48",x"c0",x"87"),
   643 => (x"f0",x"c2",x"87",x"e6"),
   644 => (x"d2",x"02",x"bf",x"d4"),
   645 => (x"c4",x"49",x"75",x"87"),
   646 => (x"cc",x"e8",x"c2",x"91"),
   647 => (x"cf",x"4c",x"69",x"81"),
   648 => (x"ff",x"ff",x"ff",x"ff"),
   649 => (x"75",x"87",x"cb",x"9c"),
   650 => (x"c2",x"91",x"c2",x"49"),
   651 => (x"9f",x"81",x"cc",x"e8"),
   652 => (x"48",x"74",x"4c",x"69"),
   653 => (x"4c",x"26",x"4d",x"26"),
   654 => (x"4f",x"26",x"4b",x"26"),
   655 => (x"5c",x"5b",x"5e",x"0e"),
   656 => (x"86",x"f4",x"0e",x"5d"),
   657 => (x"c4",x"59",x"a6",x"c8"),
   658 => (x"80",x"c8",x"48",x"66"),
   659 => (x"48",x"6e",x"7e",x"70"),
   660 => (x"c1",x"1e",x"78",x"c0"),
   661 => (x"87",x"fd",x"cc",x"49"),
   662 => (x"4c",x"70",x"86",x"c4"),
   663 => (x"fc",x"c0",x"02",x"9c"),
   664 => (x"dc",x"f0",x"c2",x"87"),
   665 => (x"49",x"66",x"dc",x"4a"),
   666 => (x"87",x"c1",x"de",x"ff"),
   667 => (x"c0",x"02",x"98",x"70"),
   668 => (x"4a",x"74",x"87",x"eb"),
   669 => (x"cb",x"49",x"66",x"dc"),
   670 => (x"cb",x"de",x"ff",x"4b"),
   671 => (x"02",x"98",x"70",x"87"),
   672 => (x"1e",x"c0",x"87",x"db"),
   673 => (x"c4",x"02",x"9c",x"74"),
   674 => (x"c2",x"4d",x"c0",x"87"),
   675 => (x"75",x"4d",x"c1",x"87"),
   676 => (x"87",x"c1",x"cc",x"49"),
   677 => (x"4c",x"70",x"86",x"c4"),
   678 => (x"c4",x"ff",x"05",x"9c"),
   679 => (x"02",x"9c",x"74",x"87"),
   680 => (x"dc",x"87",x"f4",x"c1"),
   681 => (x"48",x"6e",x"49",x"a4"),
   682 => (x"a4",x"da",x"78",x"69"),
   683 => (x"4d",x"66",x"c4",x"49"),
   684 => (x"69",x"9f",x"85",x"c4"),
   685 => (x"d4",x"f0",x"c2",x"7d"),
   686 => (x"87",x"d2",x"02",x"bf"),
   687 => (x"9f",x"49",x"a4",x"d4"),
   688 => (x"ff",x"c0",x"49",x"69"),
   689 => (x"48",x"71",x"99",x"ff"),
   690 => (x"7e",x"70",x"30",x"d0"),
   691 => (x"7e",x"c0",x"87",x"c2"),
   692 => (x"6d",x"48",x"49",x"6e"),
   693 => (x"c4",x"7d",x"70",x"80"),
   694 => (x"78",x"c0",x"48",x"66"),
   695 => (x"cc",x"49",x"66",x"c4"),
   696 => (x"c4",x"79",x"6d",x"81"),
   697 => (x"81",x"d0",x"49",x"66"),
   698 => (x"a6",x"c8",x"79",x"c0"),
   699 => (x"c8",x"78",x"c0",x"48"),
   700 => (x"66",x"c4",x"4c",x"66"),
   701 => (x"74",x"82",x"d4",x"4a"),
   702 => (x"72",x"91",x"c8",x"49"),
   703 => (x"41",x"c0",x"49",x"a1"),
   704 => (x"84",x"c1",x"79",x"6d"),
   705 => (x"04",x"ac",x"b7",x"c6"),
   706 => (x"c4",x"87",x"e7",x"ff"),
   707 => (x"c4",x"c1",x"49",x"66"),
   708 => (x"c1",x"79",x"c0",x"81"),
   709 => (x"c0",x"87",x"c2",x"48"),
   710 => (x"26",x"8e",x"f4",x"48"),
   711 => (x"26",x"4c",x"26",x"4d"),
   712 => (x"0e",x"4f",x"26",x"4b"),
   713 => (x"5d",x"5c",x"5b",x"5e"),
   714 => (x"d0",x"4c",x"71",x"0e"),
   715 => (x"49",x"6c",x"4d",x"66"),
   716 => (x"c2",x"b9",x"75",x"85"),
   717 => (x"4a",x"bf",x"d0",x"f0"),
   718 => (x"99",x"72",x"ba",x"ff"),
   719 => (x"c0",x"02",x"99",x"71"),
   720 => (x"a4",x"c4",x"87",x"e4"),
   721 => (x"f9",x"49",x"6b",x"4b"),
   722 => (x"7b",x"70",x"87",x"fb"),
   723 => (x"bf",x"cc",x"f0",x"c2"),
   724 => (x"71",x"81",x"6c",x"49"),
   725 => (x"c2",x"b9",x"75",x"7c"),
   726 => (x"4a",x"bf",x"d0",x"f0"),
   727 => (x"99",x"72",x"ba",x"ff"),
   728 => (x"ff",x"05",x"99",x"71"),
   729 => (x"7c",x"75",x"87",x"dc"),
   730 => (x"4c",x"26",x"4d",x"26"),
   731 => (x"4f",x"26",x"4b",x"26"),
   732 => (x"71",x"1e",x"73",x"1e"),
   733 => (x"f0",x"f4",x"c2",x"4b"),
   734 => (x"a3",x"c4",x"49",x"bf"),
   735 => (x"c2",x"4a",x"6a",x"4a"),
   736 => (x"cc",x"f0",x"c2",x"8a"),
   737 => (x"a1",x"72",x"92",x"bf"),
   738 => (x"d0",x"f0",x"c2",x"49"),
   739 => (x"9a",x"6b",x"4a",x"bf"),
   740 => (x"c0",x"49",x"a1",x"72"),
   741 => (x"c8",x"59",x"d4",x"fe"),
   742 => (x"e9",x"71",x"1e",x"66"),
   743 => (x"86",x"c4",x"87",x"d8"),
   744 => (x"c4",x"05",x"98",x"70"),
   745 => (x"c2",x"48",x"c0",x"87"),
   746 => (x"26",x"48",x"c1",x"87"),
   747 => (x"1e",x"4f",x"26",x"4b"),
   748 => (x"4b",x"71",x"1e",x"73"),
   749 => (x"bf",x"f0",x"f4",x"c2"),
   750 => (x"4a",x"a3",x"c4",x"49"),
   751 => (x"8a",x"c2",x"4a",x"6a"),
   752 => (x"bf",x"cc",x"f0",x"c2"),
   753 => (x"49",x"a1",x"72",x"92"),
   754 => (x"bf",x"d0",x"f0",x"c2"),
   755 => (x"72",x"9a",x"6b",x"4a"),
   756 => (x"fe",x"c0",x"49",x"a1"),
   757 => (x"66",x"c8",x"59",x"d4"),
   758 => (x"c4",x"e5",x"71",x"1e"),
   759 => (x"70",x"86",x"c4",x"87"),
   760 => (x"87",x"c4",x"05",x"98"),
   761 => (x"87",x"c2",x"48",x"c0"),
   762 => (x"4b",x"26",x"48",x"c1"),
   763 => (x"5e",x"0e",x"4f",x"26"),
   764 => (x"0e",x"5d",x"5c",x"5b"),
   765 => (x"4b",x"71",x"86",x"e4"),
   766 => (x"48",x"66",x"ec",x"c0"),
   767 => (x"a6",x"cc",x"28",x"c9"),
   768 => (x"d0",x"f0",x"c2",x"58"),
   769 => (x"b9",x"ff",x"49",x"bf"),
   770 => (x"66",x"c8",x"48",x"71"),
   771 => (x"58",x"a6",x"d4",x"98"),
   772 => (x"98",x"6b",x"48",x"71"),
   773 => (x"c4",x"58",x"a6",x"d0"),
   774 => (x"a6",x"c4",x"7e",x"a3"),
   775 => (x"78",x"bf",x"6e",x"48"),
   776 => (x"cc",x"48",x"66",x"d0"),
   777 => (x"c6",x"05",x"a8",x"66"),
   778 => (x"7b",x"66",x"c8",x"87"),
   779 => (x"d4",x"87",x"c6",x"c3"),
   780 => (x"ff",x"c1",x"48",x"a6"),
   781 => (x"ff",x"ff",x"ff",x"ff"),
   782 => (x"ff",x"80",x"c4",x"78"),
   783 => (x"d4",x"4a",x"c0",x"78"),
   784 => (x"49",x"72",x"4d",x"a3"),
   785 => (x"a1",x"75",x"91",x"c8"),
   786 => (x"4c",x"66",x"d0",x"49"),
   787 => (x"b7",x"c0",x"8c",x"69"),
   788 => (x"87",x"cd",x"04",x"ac"),
   789 => (x"ac",x"b7",x"66",x"d4"),
   790 => (x"dc",x"87",x"c6",x"03"),
   791 => (x"a6",x"d8",x"5a",x"a6"),
   792 => (x"c6",x"82",x"c1",x"5c"),
   793 => (x"ff",x"04",x"aa",x"b7"),
   794 => (x"66",x"d8",x"87",x"d5"),
   795 => (x"a8",x"b7",x"c0",x"48"),
   796 => (x"d8",x"87",x"d0",x"04"),
   797 => (x"91",x"c8",x"49",x"66"),
   798 => (x"21",x"49",x"a1",x"75"),
   799 => (x"69",x"48",x"6e",x"7b"),
   800 => (x"c0",x"87",x"c9",x"78"),
   801 => (x"49",x"a3",x"cc",x"7b"),
   802 => (x"78",x"69",x"48",x"6e"),
   803 => (x"6b",x"48",x"66",x"c8"),
   804 => (x"58",x"a6",x"cc",x"88"),
   805 => (x"bf",x"cc",x"f0",x"c2"),
   806 => (x"70",x"90",x"c8",x"48"),
   807 => (x"48",x"66",x"c8",x"7e"),
   808 => (x"c9",x"01",x"a8",x"6e"),
   809 => (x"48",x"66",x"c8",x"87"),
   810 => (x"c0",x"03",x"a8",x"6e"),
   811 => (x"c4",x"c1",x"87",x"fd"),
   812 => (x"bf",x"6e",x"7e",x"a3"),
   813 => (x"75",x"91",x"c8",x"49"),
   814 => (x"66",x"cc",x"49",x"a1"),
   815 => (x"49",x"bf",x"6e",x"79"),
   816 => (x"a1",x"75",x"91",x"c8"),
   817 => (x"66",x"81",x"c4",x"49"),
   818 => (x"48",x"a6",x"d0",x"79"),
   819 => (x"d0",x"78",x"bf",x"6e"),
   820 => (x"a8",x"c5",x"48",x"66"),
   821 => (x"c4",x"87",x"c7",x"05"),
   822 => (x"78",x"c0",x"48",x"a6"),
   823 => (x"66",x"d0",x"87",x"c8"),
   824 => (x"c8",x"80",x"c1",x"48"),
   825 => (x"48",x"6e",x"58",x"a6"),
   826 => (x"c8",x"78",x"66",x"c4"),
   827 => (x"49",x"73",x"1e",x"66"),
   828 => (x"c4",x"87",x"f0",x"f8"),
   829 => (x"cc",x"e8",x"c2",x"86"),
   830 => (x"f9",x"49",x"73",x"1e"),
   831 => (x"a3",x"d0",x"87",x"f2"),
   832 => (x"66",x"f0",x"c0",x"49"),
   833 => (x"26",x"8e",x"e0",x"79"),
   834 => (x"26",x"4c",x"26",x"4d"),
   835 => (x"0e",x"4f",x"26",x"4b"),
   836 => (x"0e",x"5c",x"5b",x"5e"),
   837 => (x"4b",x"c0",x"4a",x"71"),
   838 => (x"c0",x"02",x"9a",x"72"),
   839 => (x"a2",x"da",x"87",x"e0"),
   840 => (x"4b",x"69",x"9f",x"49"),
   841 => (x"bf",x"d4",x"f0",x"c2"),
   842 => (x"d4",x"87",x"cf",x"02"),
   843 => (x"69",x"9f",x"49",x"a2"),
   844 => (x"ff",x"c0",x"4c",x"49"),
   845 => (x"34",x"d0",x"9c",x"ff"),
   846 => (x"4c",x"c0",x"87",x"c2"),
   847 => (x"9b",x"73",x"b3",x"74"),
   848 => (x"4a",x"87",x"df",x"02"),
   849 => (x"f0",x"c2",x"8a",x"c2"),
   850 => (x"92",x"49",x"bf",x"cc"),
   851 => (x"bf",x"f0",x"f4",x"c2"),
   852 => (x"c2",x"80",x"72",x"48"),
   853 => (x"71",x"58",x"d0",x"f5"),
   854 => (x"c2",x"30",x"c4",x"48"),
   855 => (x"c0",x"58",x"dc",x"f0"),
   856 => (x"f4",x"c2",x"87",x"e9"),
   857 => (x"c2",x"4b",x"bf",x"f4"),
   858 => (x"c2",x"48",x"cc",x"f5"),
   859 => (x"78",x"bf",x"f8",x"f4"),
   860 => (x"bf",x"d4",x"f0",x"c2"),
   861 => (x"c2",x"87",x"c9",x"02"),
   862 => (x"49",x"bf",x"cc",x"f0"),
   863 => (x"87",x"c7",x"31",x"c4"),
   864 => (x"bf",x"fc",x"f4",x"c2"),
   865 => (x"c2",x"31",x"c4",x"49"),
   866 => (x"c2",x"59",x"dc",x"f0"),
   867 => (x"26",x"5b",x"cc",x"f5"),
   868 => (x"26",x"4b",x"26",x"4c"),
   869 => (x"5b",x"5e",x"0e",x"4f"),
   870 => (x"f0",x"0e",x"5d",x"5c"),
   871 => (x"59",x"a6",x"c8",x"86"),
   872 => (x"ff",x"ff",x"ff",x"cf"),
   873 => (x"7e",x"c0",x"4c",x"f8"),
   874 => (x"d8",x"02",x"66",x"c4"),
   875 => (x"c8",x"e8",x"c2",x"87"),
   876 => (x"c2",x"78",x"c0",x"48"),
   877 => (x"c2",x"48",x"c0",x"e8"),
   878 => (x"78",x"bf",x"cc",x"f5"),
   879 => (x"48",x"c4",x"e8",x"c2"),
   880 => (x"bf",x"c8",x"f5",x"c2"),
   881 => (x"e9",x"f0",x"c2",x"78"),
   882 => (x"c2",x"50",x"c0",x"48"),
   883 => (x"49",x"bf",x"d8",x"f0"),
   884 => (x"bf",x"c8",x"e8",x"c2"),
   885 => (x"03",x"aa",x"71",x"4a"),
   886 => (x"72",x"87",x"cc",x"c4"),
   887 => (x"05",x"99",x"cf",x"49"),
   888 => (x"c0",x"87",x"ea",x"c0"),
   889 => (x"c2",x"48",x"d0",x"fe"),
   890 => (x"78",x"bf",x"c0",x"e8"),
   891 => (x"1e",x"cc",x"e8",x"c2"),
   892 => (x"bf",x"c0",x"e8",x"c2"),
   893 => (x"c0",x"e8",x"c2",x"49"),
   894 => (x"78",x"a1",x"c1",x"48"),
   895 => (x"f5",x"df",x"ff",x"71"),
   896 => (x"c0",x"86",x"c4",x"87"),
   897 => (x"c2",x"48",x"cc",x"fe"),
   898 => (x"cc",x"78",x"cc",x"e8"),
   899 => (x"cc",x"fe",x"c0",x"87"),
   900 => (x"e0",x"c0",x"48",x"bf"),
   901 => (x"d0",x"fe",x"c0",x"80"),
   902 => (x"c8",x"e8",x"c2",x"58"),
   903 => (x"80",x"c1",x"48",x"bf"),
   904 => (x"58",x"cc",x"e8",x"c2"),
   905 => (x"00",x"0f",x"8c",x"27"),
   906 => (x"bf",x"97",x"bf",x"00"),
   907 => (x"c2",x"02",x"9d",x"4d"),
   908 => (x"e5",x"c3",x"87",x"e5"),
   909 => (x"de",x"c2",x"02",x"ad"),
   910 => (x"cc",x"fe",x"c0",x"87"),
   911 => (x"a3",x"cb",x"4b",x"bf"),
   912 => (x"cf",x"4c",x"11",x"49"),
   913 => (x"d2",x"c1",x"05",x"ac"),
   914 => (x"df",x"49",x"75",x"87"),
   915 => (x"cd",x"89",x"c1",x"99"),
   916 => (x"dc",x"f0",x"c2",x"91"),
   917 => (x"4a",x"a3",x"c1",x"81"),
   918 => (x"a3",x"c3",x"51",x"12"),
   919 => (x"c5",x"51",x"12",x"4a"),
   920 => (x"51",x"12",x"4a",x"a3"),
   921 => (x"12",x"4a",x"a3",x"c7"),
   922 => (x"4a",x"a3",x"c9",x"51"),
   923 => (x"a3",x"ce",x"51",x"12"),
   924 => (x"d0",x"51",x"12",x"4a"),
   925 => (x"51",x"12",x"4a",x"a3"),
   926 => (x"12",x"4a",x"a3",x"d2"),
   927 => (x"4a",x"a3",x"d4",x"51"),
   928 => (x"a3",x"d6",x"51",x"12"),
   929 => (x"d8",x"51",x"12",x"4a"),
   930 => (x"51",x"12",x"4a",x"a3"),
   931 => (x"12",x"4a",x"a3",x"dc"),
   932 => (x"4a",x"a3",x"de",x"51"),
   933 => (x"7e",x"c1",x"51",x"12"),
   934 => (x"74",x"87",x"fc",x"c0"),
   935 => (x"05",x"99",x"c8",x"49"),
   936 => (x"74",x"87",x"ed",x"c0"),
   937 => (x"05",x"99",x"d0",x"49"),
   938 => (x"e0",x"c0",x"87",x"d3"),
   939 => (x"cc",x"c0",x"02",x"66"),
   940 => (x"c0",x"49",x"73",x"87"),
   941 => (x"70",x"0f",x"66",x"e0"),
   942 => (x"d3",x"c0",x"02",x"98"),
   943 => (x"c0",x"05",x"6e",x"87"),
   944 => (x"f0",x"c2",x"87",x"c6"),
   945 => (x"50",x"c0",x"48",x"dc"),
   946 => (x"bf",x"cc",x"fe",x"c0"),
   947 => (x"87",x"e9",x"c2",x"48"),
   948 => (x"48",x"e9",x"f0",x"c2"),
   949 => (x"c2",x"7e",x"50",x"c0"),
   950 => (x"49",x"bf",x"d8",x"f0"),
   951 => (x"bf",x"c8",x"e8",x"c2"),
   952 => (x"04",x"aa",x"71",x"4a"),
   953 => (x"cf",x"87",x"f4",x"fb"),
   954 => (x"f8",x"ff",x"ff",x"ff"),
   955 => (x"cc",x"f5",x"c2",x"4c"),
   956 => (x"c8",x"c0",x"05",x"bf"),
   957 => (x"d4",x"f0",x"c2",x"87"),
   958 => (x"fa",x"c1",x"02",x"bf"),
   959 => (x"c4",x"e8",x"c2",x"87"),
   960 => (x"c0",x"eb",x"49",x"bf"),
   961 => (x"c8",x"e8",x"c2",x"87"),
   962 => (x"48",x"a6",x"c4",x"58"),
   963 => (x"bf",x"c4",x"e8",x"c2"),
   964 => (x"d4",x"f0",x"c2",x"78"),
   965 => (x"db",x"c0",x"02",x"bf"),
   966 => (x"49",x"66",x"c4",x"87"),
   967 => (x"a9",x"74",x"99",x"74"),
   968 => (x"87",x"c8",x"c0",x"02"),
   969 => (x"c0",x"48",x"a6",x"c8"),
   970 => (x"87",x"e7",x"c0",x"78"),
   971 => (x"c1",x"48",x"a6",x"c8"),
   972 => (x"87",x"df",x"c0",x"78"),
   973 => (x"cf",x"49",x"66",x"c4"),
   974 => (x"a9",x"99",x"f8",x"ff"),
   975 => (x"87",x"c8",x"c0",x"02"),
   976 => (x"c0",x"48",x"a6",x"cc"),
   977 => (x"87",x"c5",x"c0",x"78"),
   978 => (x"c1",x"48",x"a6",x"cc"),
   979 => (x"48",x"a6",x"c8",x"78"),
   980 => (x"c8",x"78",x"66",x"cc"),
   981 => (x"de",x"c0",x"05",x"66"),
   982 => (x"49",x"66",x"c4",x"87"),
   983 => (x"f0",x"c2",x"89",x"c2"),
   984 => (x"c2",x"91",x"bf",x"cc"),
   985 => (x"48",x"bf",x"f0",x"f4"),
   986 => (x"e8",x"c2",x"80",x"71"),
   987 => (x"e8",x"c2",x"58",x"c4"),
   988 => (x"78",x"c0",x"48",x"c8"),
   989 => (x"c0",x"87",x"d4",x"f9"),
   990 => (x"ff",x"ff",x"cf",x"48"),
   991 => (x"f0",x"4c",x"f8",x"ff"),
   992 => (x"26",x"4d",x"26",x"8e"),
   993 => (x"26",x"4b",x"26",x"4c"),
   994 => (x"00",x"00",x"00",x"4f"),
   995 => (x"00",x"00",x"00",x"00"),
   996 => (x"ff",x"ff",x"ff",x"ff"),
   997 => (x"48",x"d4",x"ff",x"1e"),
   998 => (x"68",x"78",x"ff",x"c3"),
   999 => (x"1e",x"4f",x"26",x"48"),
  1000 => (x"c3",x"48",x"d4",x"ff"),
  1001 => (x"d0",x"ff",x"78",x"ff"),
  1002 => (x"78",x"e1",x"c0",x"48"),
  1003 => (x"d4",x"48",x"d4",x"ff"),
  1004 => (x"1e",x"4f",x"26",x"78"),
  1005 => (x"c0",x"48",x"d0",x"ff"),
  1006 => (x"4f",x"26",x"78",x"e0"),
  1007 => (x"87",x"d4",x"ff",x"1e"),
  1008 => (x"02",x"99",x"49",x"70"),
  1009 => (x"fb",x"c0",x"87",x"c6"),
  1010 => (x"87",x"f1",x"05",x"a9"),
  1011 => (x"4f",x"26",x"48",x"71"),
  1012 => (x"5c",x"5b",x"5e",x"0e"),
  1013 => (x"c0",x"4b",x"71",x"0e"),
  1014 => (x"87",x"f8",x"fe",x"4c"),
  1015 => (x"02",x"99",x"49",x"70"),
  1016 => (x"c0",x"87",x"f9",x"c0"),
  1017 => (x"c0",x"02",x"a9",x"ec"),
  1018 => (x"fb",x"c0",x"87",x"f2"),
  1019 => (x"eb",x"c0",x"02",x"a9"),
  1020 => (x"b7",x"66",x"cc",x"87"),
  1021 => (x"87",x"c7",x"03",x"ac"),
  1022 => (x"c2",x"02",x"66",x"d0"),
  1023 => (x"71",x"53",x"71",x"87"),
  1024 => (x"87",x"c2",x"02",x"99"),
  1025 => (x"cb",x"fe",x"84",x"c1"),
  1026 => (x"99",x"49",x"70",x"87"),
  1027 => (x"c0",x"87",x"cd",x"02"),
  1028 => (x"c7",x"02",x"a9",x"ec"),
  1029 => (x"a9",x"fb",x"c0",x"87"),
  1030 => (x"87",x"d5",x"ff",x"05"),
  1031 => (x"c3",x"02",x"66",x"d0"),
  1032 => (x"7b",x"97",x"c0",x"87"),
  1033 => (x"05",x"a9",x"fb",x"c0"),
  1034 => (x"4a",x"74",x"87",x"c7"),
  1035 => (x"c2",x"8a",x"0a",x"c0"),
  1036 => (x"72",x"4a",x"74",x"87"),
  1037 => (x"26",x"4c",x"26",x"48"),
  1038 => (x"1e",x"4f",x"26",x"4b"),
  1039 => (x"70",x"87",x"d5",x"fd"),
  1040 => (x"a9",x"f0",x"c0",x"49"),
  1041 => (x"c0",x"87",x"c9",x"04"),
  1042 => (x"c3",x"01",x"a9",x"f9"),
  1043 => (x"89",x"f0",x"c0",x"87"),
  1044 => (x"04",x"a9",x"c1",x"c1"),
  1045 => (x"da",x"c1",x"87",x"c9"),
  1046 => (x"87",x"c3",x"01",x"a9"),
  1047 => (x"71",x"89",x"f7",x"c0"),
  1048 => (x"0e",x"4f",x"26",x"48"),
  1049 => (x"5d",x"5c",x"5b",x"5e"),
  1050 => (x"71",x"86",x"f8",x"0e"),
  1051 => (x"fc",x"7e",x"c0",x"4c"),
  1052 => (x"4b",x"c0",x"87",x"ed"),
  1053 => (x"97",x"c4",x"c4",x"c1"),
  1054 => (x"a9",x"c0",x"49",x"bf"),
  1055 => (x"fc",x"87",x"cf",x"04"),
  1056 => (x"83",x"c1",x"87",x"fa"),
  1057 => (x"97",x"c4",x"c4",x"c1"),
  1058 => (x"06",x"ab",x"49",x"bf"),
  1059 => (x"c4",x"c1",x"87",x"f1"),
  1060 => (x"02",x"bf",x"97",x"c4"),
  1061 => (x"fb",x"fb",x"87",x"cf"),
  1062 => (x"99",x"49",x"70",x"87"),
  1063 => (x"c0",x"87",x"c6",x"02"),
  1064 => (x"f1",x"05",x"a9",x"ec"),
  1065 => (x"fb",x"4b",x"c0",x"87"),
  1066 => (x"4d",x"70",x"87",x"ea"),
  1067 => (x"c8",x"87",x"e5",x"fb"),
  1068 => (x"df",x"fb",x"58",x"a6"),
  1069 => (x"c1",x"4a",x"70",x"87"),
  1070 => (x"49",x"a4",x"c8",x"83"),
  1071 => (x"ad",x"49",x"69",x"97"),
  1072 => (x"c9",x"87",x"da",x"05"),
  1073 => (x"69",x"97",x"49",x"a4"),
  1074 => (x"a9",x"66",x"c4",x"49"),
  1075 => (x"ca",x"87",x"ce",x"05"),
  1076 => (x"69",x"97",x"49",x"a4"),
  1077 => (x"c4",x"05",x"aa",x"49"),
  1078 => (x"d0",x"7e",x"c1",x"87"),
  1079 => (x"ad",x"ec",x"c0",x"87"),
  1080 => (x"c0",x"87",x"c6",x"02"),
  1081 => (x"c4",x"05",x"ad",x"fb"),
  1082 => (x"c1",x"4b",x"c0",x"87"),
  1083 => (x"fe",x"02",x"6e",x"7e"),
  1084 => (x"fe",x"fa",x"87",x"f5"),
  1085 => (x"f8",x"48",x"73",x"87"),
  1086 => (x"26",x"4d",x"26",x"8e"),
  1087 => (x"26",x"4b",x"26",x"4c"),
  1088 => (x"00",x"00",x"00",x"4f"),
  1089 => (x"1e",x"73",x"1e",x"00"),
  1090 => (x"c8",x"4b",x"d4",x"ff"),
  1091 => (x"d0",x"ff",x"4a",x"66"),
  1092 => (x"78",x"c5",x"c8",x"48"),
  1093 => (x"c1",x"48",x"d4",x"ff"),
  1094 => (x"7b",x"11",x"78",x"d4"),
  1095 => (x"f9",x"05",x"8a",x"c1"),
  1096 => (x"48",x"d0",x"ff",x"87"),
  1097 => (x"4b",x"26",x"78",x"c4"),
  1098 => (x"5e",x"0e",x"4f",x"26"),
  1099 => (x"0e",x"5d",x"5c",x"5b"),
  1100 => (x"7e",x"71",x"86",x"f8"),
  1101 => (x"f5",x"c2",x"1e",x"6e"),
  1102 => (x"ff",x"e3",x"49",x"e0"),
  1103 => (x"70",x"86",x"c4",x"87"),
  1104 => (x"ed",x"c4",x"02",x"98"),
  1105 => (x"f4",x"f1",x"c1",x"87"),
  1106 => (x"49",x"6e",x"4c",x"bf"),
  1107 => (x"c8",x"87",x"d4",x"fc"),
  1108 => (x"ca",x"c1",x"58",x"a6"),
  1109 => (x"fc",x"fe",x"1e",x"c0"),
  1110 => (x"86",x"c4",x"87",x"f2"),
  1111 => (x"87",x"c5",x"05",x"66"),
  1112 => (x"c1",x"48",x"a6",x"c4"),
  1113 => (x"48",x"d0",x"ff",x"78"),
  1114 => (x"d4",x"ff",x"78",x"c5"),
  1115 => (x"78",x"d5",x"c1",x"48"),
  1116 => (x"c1",x"49",x"66",x"c4"),
  1117 => (x"c1",x"31",x"c6",x"89"),
  1118 => (x"bf",x"97",x"ec",x"f1"),
  1119 => (x"b0",x"71",x"48",x"4a"),
  1120 => (x"78",x"08",x"d4",x"ff"),
  1121 => (x"c4",x"48",x"d0",x"ff"),
  1122 => (x"dc",x"f5",x"c2",x"78"),
  1123 => (x"d0",x"49",x"bf",x"97"),
  1124 => (x"87",x"dd",x"02",x"99"),
  1125 => (x"d4",x"ff",x"78",x"c5"),
  1126 => (x"78",x"d6",x"c1",x"48"),
  1127 => (x"d4",x"ff",x"4a",x"c0"),
  1128 => (x"78",x"ff",x"c3",x"48"),
  1129 => (x"e0",x"c0",x"82",x"c1"),
  1130 => (x"87",x"f2",x"04",x"aa"),
  1131 => (x"c4",x"48",x"d0",x"ff"),
  1132 => (x"48",x"d4",x"ff",x"78"),
  1133 => (x"ff",x"78",x"ff",x"c3"),
  1134 => (x"78",x"c5",x"48",x"d0"),
  1135 => (x"c1",x"48",x"d4",x"ff"),
  1136 => (x"78",x"c1",x"78",x"d3"),
  1137 => (x"c4",x"48",x"d0",x"ff"),
  1138 => (x"ac",x"b7",x"c0",x"78"),
  1139 => (x"87",x"cb",x"c2",x"06"),
  1140 => (x"bf",x"e8",x"f5",x"c2"),
  1141 => (x"7e",x"74",x"8c",x"4b"),
  1142 => (x"c1",x"02",x"9b",x"73"),
  1143 => (x"c0",x"c8",x"87",x"dd"),
  1144 => (x"b7",x"c0",x"8b",x"4d"),
  1145 => (x"87",x"c6",x"03",x"ab"),
  1146 => (x"4d",x"a3",x"c0",x"c8"),
  1147 => (x"f5",x"c2",x"4b",x"c0"),
  1148 => (x"49",x"bf",x"97",x"dc"),
  1149 => (x"cf",x"02",x"99",x"d0"),
  1150 => (x"c2",x"1e",x"c0",x"87"),
  1151 => (x"e5",x"49",x"e0",x"f5"),
  1152 => (x"86",x"c4",x"87",x"ee"),
  1153 => (x"87",x"d8",x"4c",x"70"),
  1154 => (x"1e",x"cc",x"e8",x"c2"),
  1155 => (x"49",x"e0",x"f5",x"c2"),
  1156 => (x"70",x"87",x"dd",x"e5"),
  1157 => (x"c2",x"1e",x"75",x"4c"),
  1158 => (x"fb",x"49",x"cc",x"e8"),
  1159 => (x"86",x"c8",x"87",x"e7"),
  1160 => (x"c5",x"05",x"9c",x"74"),
  1161 => (x"c1",x"48",x"c0",x"87"),
  1162 => (x"1e",x"c1",x"87",x"ca"),
  1163 => (x"49",x"e0",x"f5",x"c2"),
  1164 => (x"c4",x"87",x"f0",x"e3"),
  1165 => (x"05",x"9b",x"73",x"86"),
  1166 => (x"6e",x"87",x"e3",x"fe"),
  1167 => (x"ac",x"b7",x"c0",x"4c"),
  1168 => (x"c2",x"87",x"d1",x"06"),
  1169 => (x"c0",x"48",x"e0",x"f5"),
  1170 => (x"c0",x"80",x"d0",x"78"),
  1171 => (x"c2",x"80",x"f4",x"78"),
  1172 => (x"78",x"bf",x"ec",x"f5"),
  1173 => (x"01",x"ac",x"b7",x"c0"),
  1174 => (x"ff",x"87",x"f5",x"fd"),
  1175 => (x"78",x"c5",x"48",x"d0"),
  1176 => (x"c1",x"48",x"d4",x"ff"),
  1177 => (x"78",x"c0",x"78",x"d3"),
  1178 => (x"c4",x"48",x"d0",x"ff"),
  1179 => (x"c0",x"48",x"c1",x"78"),
  1180 => (x"48",x"c0",x"87",x"c2"),
  1181 => (x"4d",x"26",x"8e",x"f8"),
  1182 => (x"4b",x"26",x"4c",x"26"),
  1183 => (x"00",x"00",x"4f",x"26"),
  1184 => (x"20",x"74",x"6f",x"47"),
  1185 => (x"69",x"74",x"78",x"65"),
  1186 => (x"00",x"00",x"64",x"6e"),
  1187 => (x"64",x"61",x"6f",x"4c"),
  1188 => (x"2e",x"67",x"6e",x"69"),
  1189 => (x"00",x"00",x"2e",x"2e"),
  1190 => (x"61",x"42",x"20",x"80"),
  1191 => (x"00",x"00",x"6b",x"63"),
  1192 => (x"64",x"61",x"6f",x"4c"),
  1193 => (x"20",x"2e",x"2a",x"20"),
  1194 => (x"00",x"00",x"00",x"00"),
  1195 => (x"00",x"00",x"20",x"3a"),
  1196 => (x"61",x"42",x"20",x"80"),
  1197 => (x"00",x"00",x"6b",x"63"),
  1198 => (x"78",x"45",x"20",x"80"),
  1199 => (x"00",x"00",x"74",x"69"),
  1200 => (x"49",x"20",x"44",x"53"),
  1201 => (x"2e",x"74",x"69",x"6e"),
  1202 => (x"00",x"00",x"00",x"2e"),
  1203 => (x"00",x"00",x"4b",x"4f"),
  1204 => (x"54",x"4f",x"4f",x"42"),
  1205 => (x"20",x"20",x"20",x"20"),
  1206 => (x"00",x"4d",x"4f",x"52"),
  1207 => (x"5c",x"5b",x"5e",x"0e"),
  1208 => (x"86",x"fc",x"0e",x"5d"),
  1209 => (x"4b",x"c0",x"4d",x"71"),
  1210 => (x"c0",x"04",x"ad",x"4c"),
  1211 => (x"c1",x"c1",x"87",x"e8"),
  1212 => (x"9c",x"74",x"1e",x"e3"),
  1213 => (x"c0",x"87",x"c4",x"02"),
  1214 => (x"c1",x"87",x"c2",x"4a"),
  1215 => (x"ea",x"49",x"72",x"4a"),
  1216 => (x"86",x"c4",x"87",x"d3"),
  1217 => (x"83",x"c1",x"7e",x"70"),
  1218 => (x"87",x"c2",x"05",x"6e"),
  1219 => (x"84",x"c1",x"4b",x"75"),
  1220 => (x"ff",x"06",x"ab",x"75"),
  1221 => (x"48",x"6e",x"87",x"d8"),
  1222 => (x"4d",x"26",x"8e",x"fc"),
  1223 => (x"4b",x"26",x"4c",x"26"),
  1224 => (x"5e",x"0e",x"4f",x"26"),
  1225 => (x"71",x"0e",x"5c",x"5b"),
  1226 => (x"02",x"66",x"cc",x"4b"),
  1227 => (x"c0",x"4c",x"87",x"d8"),
  1228 => (x"d8",x"02",x"8c",x"f0"),
  1229 => (x"c1",x"4a",x"74",x"87"),
  1230 => (x"87",x"d1",x"02",x"8a"),
  1231 => (x"87",x"cd",x"02",x"8a"),
  1232 => (x"87",x"c9",x"02",x"8a"),
  1233 => (x"49",x"73",x"87",x"d9"),
  1234 => (x"d2",x"87",x"df",x"f7"),
  1235 => (x"c0",x"1e",x"74",x"87"),
  1236 => (x"db",x"d7",x"c1",x"49"),
  1237 => (x"73",x"1e",x"74",x"87"),
  1238 => (x"d3",x"d7",x"c1",x"49"),
  1239 => (x"26",x"86",x"c8",x"87"),
  1240 => (x"26",x"4b",x"26",x"4c"),
  1241 => (x"5b",x"5e",x"0e",x"4f"),
  1242 => (x"fc",x"0e",x"5d",x"5c"),
  1243 => (x"49",x"4c",x"71",x"86"),
  1244 => (x"f7",x"c2",x"91",x"de"),
  1245 => (x"85",x"71",x"4d",x"c0"),
  1246 => (x"c1",x"02",x"6d",x"97"),
  1247 => (x"f6",x"c2",x"87",x"db"),
  1248 => (x"74",x"49",x"bf",x"f0"),
  1249 => (x"d3",x"fd",x"71",x"81"),
  1250 => (x"48",x"7e",x"70",x"87"),
  1251 => (x"f2",x"c0",x"02",x"98"),
  1252 => (x"f4",x"f6",x"c2",x"87"),
  1253 => (x"cb",x"4a",x"70",x"4b"),
  1254 => (x"c5",x"fa",x"fe",x"49"),
  1255 => (x"cc",x"4b",x"74",x"87"),
  1256 => (x"f8",x"f1",x"c1",x"93"),
  1257 => (x"c1",x"83",x"c4",x"83"),
  1258 => (x"74",x"7b",x"cc",x"ca"),
  1259 => (x"cb",x"c1",x"c1",x"49"),
  1260 => (x"c1",x"7b",x"75",x"87"),
  1261 => (x"bf",x"97",x"f0",x"f1"),
  1262 => (x"f6",x"c2",x"1e",x"49"),
  1263 => (x"e1",x"fd",x"49",x"f4"),
  1264 => (x"74",x"86",x"c4",x"87"),
  1265 => (x"f3",x"c0",x"c1",x"49"),
  1266 => (x"c1",x"49",x"c0",x"87"),
  1267 => (x"c2",x"87",x"ce",x"c2"),
  1268 => (x"c0",x"48",x"d8",x"f5"),
  1269 => (x"e4",x"df",x"49",x"50"),
  1270 => (x"26",x"8e",x"fc",x"87"),
  1271 => (x"26",x"4c",x"26",x"4d"),
  1272 => (x"1e",x"4f",x"26",x"4b"),
  1273 => (x"4b",x"71",x"1e",x"73"),
  1274 => (x"f0",x"f6",x"c2",x"49"),
  1275 => (x"fb",x"71",x"81",x"bf"),
  1276 => (x"4a",x"70",x"87",x"ea"),
  1277 => (x"87",x"c4",x"02",x"9a"),
  1278 => (x"87",x"d3",x"e4",x"49"),
  1279 => (x"48",x"f0",x"f6",x"c2"),
  1280 => (x"49",x"73",x"78",x"c0"),
  1281 => (x"26",x"87",x"fa",x"c1"),
  1282 => (x"1e",x"4f",x"26",x"4b"),
  1283 => (x"4b",x"71",x"1e",x"73"),
  1284 => (x"02",x"4a",x"a3",x"c4"),
  1285 => (x"c1",x"87",x"d0",x"c1"),
  1286 => (x"87",x"dc",x"02",x"8a"),
  1287 => (x"f2",x"c0",x"02",x"8a"),
  1288 => (x"c1",x"05",x"8a",x"87"),
  1289 => (x"f6",x"c2",x"87",x"d3"),
  1290 => (x"c1",x"02",x"bf",x"f0"),
  1291 => (x"c1",x"48",x"87",x"cb"),
  1292 => (x"f4",x"f6",x"c2",x"88"),
  1293 => (x"87",x"c1",x"c1",x"58"),
  1294 => (x"bf",x"f0",x"f6",x"c2"),
  1295 => (x"c2",x"89",x"c6",x"49"),
  1296 => (x"c0",x"59",x"f4",x"f6"),
  1297 => (x"c0",x"03",x"a9",x"b7"),
  1298 => (x"f6",x"c2",x"87",x"ef"),
  1299 => (x"78",x"c0",x"48",x"f0"),
  1300 => (x"c2",x"87",x"e6",x"c0"),
  1301 => (x"02",x"bf",x"ec",x"f6"),
  1302 => (x"f6",x"c2",x"87",x"df"),
  1303 => (x"c1",x"48",x"bf",x"f0"),
  1304 => (x"f4",x"f6",x"c2",x"80"),
  1305 => (x"c2",x"87",x"d2",x"58"),
  1306 => (x"02",x"bf",x"ec",x"f6"),
  1307 => (x"f6",x"c2",x"87",x"cb"),
  1308 => (x"c6",x"48",x"bf",x"f0"),
  1309 => (x"f4",x"f6",x"c2",x"80"),
  1310 => (x"c4",x"49",x"73",x"58"),
  1311 => (x"26",x"4b",x"26",x"87"),
  1312 => (x"5b",x"5e",x"0e",x"4f"),
  1313 => (x"f0",x"0e",x"5d",x"5c"),
  1314 => (x"59",x"a6",x"d0",x"86"),
  1315 => (x"4d",x"cc",x"e8",x"c2"),
  1316 => (x"f6",x"c2",x"4c",x"c0"),
  1317 => (x"78",x"c1",x"48",x"ec"),
  1318 => (x"c0",x"48",x"a6",x"c8"),
  1319 => (x"c2",x"7e",x"75",x"78"),
  1320 => (x"48",x"bf",x"f0",x"f6"),
  1321 => (x"c1",x"06",x"a8",x"c0"),
  1322 => (x"a6",x"c8",x"87",x"c0"),
  1323 => (x"c2",x"7e",x"75",x"5c"),
  1324 => (x"98",x"48",x"cc",x"e8"),
  1325 => (x"87",x"f2",x"c0",x"02"),
  1326 => (x"c1",x"4d",x"66",x"c4"),
  1327 => (x"cc",x"1e",x"e3",x"c1"),
  1328 => (x"87",x"c4",x"02",x"66"),
  1329 => (x"87",x"c2",x"4c",x"c0"),
  1330 => (x"49",x"74",x"4c",x"c1"),
  1331 => (x"c4",x"87",x"c6",x"e3"),
  1332 => (x"c1",x"7e",x"70",x"86"),
  1333 => (x"48",x"66",x"c8",x"85"),
  1334 => (x"a6",x"cc",x"80",x"c1"),
  1335 => (x"f0",x"f6",x"c2",x"58"),
  1336 => (x"c5",x"03",x"ad",x"bf"),
  1337 => (x"ff",x"05",x"6e",x"87"),
  1338 => (x"4d",x"6e",x"87",x"d1"),
  1339 => (x"9d",x"75",x"4c",x"c0"),
  1340 => (x"87",x"dc",x"c3",x"02"),
  1341 => (x"1e",x"e3",x"c1",x"c1"),
  1342 => (x"c7",x"02",x"66",x"cc"),
  1343 => (x"48",x"a6",x"c8",x"87"),
  1344 => (x"87",x"c5",x"78",x"c0"),
  1345 => (x"c1",x"48",x"a6",x"c8"),
  1346 => (x"49",x"66",x"c8",x"78"),
  1347 => (x"c4",x"87",x"c6",x"e2"),
  1348 => (x"48",x"7e",x"70",x"86"),
  1349 => (x"e4",x"c2",x"02",x"98"),
  1350 => (x"81",x"cb",x"49",x"87"),
  1351 => (x"d0",x"49",x"69",x"97"),
  1352 => (x"d4",x"c1",x"02",x"99"),
  1353 => (x"cc",x"49",x"74",x"87"),
  1354 => (x"f8",x"f1",x"c1",x"91"),
  1355 => (x"e3",x"cf",x"c1",x"81"),
  1356 => (x"c3",x"81",x"c8",x"79"),
  1357 => (x"49",x"74",x"51",x"ff"),
  1358 => (x"f7",x"c2",x"91",x"de"),
  1359 => (x"85",x"71",x"4d",x"c0"),
  1360 => (x"7d",x"97",x"c1",x"c2"),
  1361 => (x"c0",x"49",x"a5",x"c1"),
  1362 => (x"f0",x"c2",x"51",x"e0"),
  1363 => (x"02",x"bf",x"97",x"dc"),
  1364 => (x"84",x"c1",x"87",x"d2"),
  1365 => (x"c2",x"4b",x"a5",x"c2"),
  1366 => (x"db",x"4a",x"dc",x"f0"),
  1367 => (x"c1",x"f3",x"fe",x"49"),
  1368 => (x"87",x"d9",x"c1",x"87"),
  1369 => (x"c0",x"49",x"a5",x"cd"),
  1370 => (x"c2",x"84",x"c1",x"51"),
  1371 => (x"4a",x"6e",x"4b",x"a5"),
  1372 => (x"f2",x"fe",x"49",x"cb"),
  1373 => (x"c4",x"c1",x"87",x"ec"),
  1374 => (x"cc",x"49",x"74",x"87"),
  1375 => (x"f8",x"f1",x"c1",x"91"),
  1376 => (x"e5",x"cd",x"c1",x"81"),
  1377 => (x"dc",x"f0",x"c2",x"79"),
  1378 => (x"d8",x"02",x"bf",x"97"),
  1379 => (x"de",x"49",x"74",x"87"),
  1380 => (x"c2",x"84",x"c1",x"91"),
  1381 => (x"71",x"4b",x"c0",x"f7"),
  1382 => (x"dc",x"f0",x"c2",x"83"),
  1383 => (x"fe",x"49",x"dd",x"4a"),
  1384 => (x"d8",x"87",x"ff",x"f1"),
  1385 => (x"de",x"4b",x"74",x"87"),
  1386 => (x"c0",x"f7",x"c2",x"93"),
  1387 => (x"49",x"a3",x"cb",x"83"),
  1388 => (x"84",x"c1",x"51",x"c0"),
  1389 => (x"cb",x"4a",x"6e",x"73"),
  1390 => (x"e5",x"f1",x"fe",x"49"),
  1391 => (x"48",x"66",x"c8",x"87"),
  1392 => (x"a6",x"cc",x"80",x"c1"),
  1393 => (x"03",x"ac",x"c7",x"58"),
  1394 => (x"6e",x"87",x"c5",x"c0"),
  1395 => (x"87",x"e4",x"fc",x"05"),
  1396 => (x"c0",x"03",x"ac",x"c7"),
  1397 => (x"f6",x"c2",x"87",x"e4"),
  1398 => (x"78",x"c0",x"48",x"ec"),
  1399 => (x"91",x"cc",x"49",x"74"),
  1400 => (x"81",x"f8",x"f1",x"c1"),
  1401 => (x"79",x"e5",x"cd",x"c1"),
  1402 => (x"91",x"de",x"49",x"74"),
  1403 => (x"81",x"c0",x"f7",x"c2"),
  1404 => (x"84",x"c1",x"51",x"c0"),
  1405 => (x"ff",x"04",x"ac",x"c7"),
  1406 => (x"f3",x"c1",x"87",x"dc"),
  1407 => (x"50",x"c0",x"48",x"d4"),
  1408 => (x"d9",x"c1",x"80",x"f7"),
  1409 => (x"ca",x"c1",x"40",x"d9"),
  1410 => (x"80",x"c8",x"78",x"d8"),
  1411 => (x"78",x"cb",x"d0",x"c1"),
  1412 => (x"c0",x"49",x"66",x"cc"),
  1413 => (x"f0",x"87",x"e5",x"f7"),
  1414 => (x"26",x"4d",x"26",x"8e"),
  1415 => (x"26",x"4b",x"26",x"4c"),
  1416 => (x"1e",x"73",x"1e",x"4f"),
  1417 => (x"cc",x"49",x"4b",x"71"),
  1418 => (x"f8",x"f1",x"c1",x"91"),
  1419 => (x"4a",x"a1",x"c8",x"81"),
  1420 => (x"48",x"ec",x"f1",x"c1"),
  1421 => (x"a1",x"c9",x"50",x"12"),
  1422 => (x"c4",x"c4",x"c1",x"4a"),
  1423 => (x"ca",x"50",x"12",x"48"),
  1424 => (x"f0",x"f1",x"c1",x"81"),
  1425 => (x"73",x"50",x"11",x"48"),
  1426 => (x"87",x"f5",x"f8",x"49"),
  1427 => (x"4f",x"26",x"4b",x"26"),
  1428 => (x"c0",x"49",x"c0",x"1e"),
  1429 => (x"26",x"87",x"c6",x"f8"),
  1430 => (x"4a",x"71",x"1e",x"4f"),
  1431 => (x"c1",x"91",x"cc",x"49"),
  1432 => (x"c8",x"81",x"f8",x"f1"),
  1433 => (x"d8",x"f5",x"c2",x"81"),
  1434 => (x"c0",x"50",x"11",x"48"),
  1435 => (x"fe",x"49",x"a2",x"f0"),
  1436 => (x"c0",x"87",x"fb",x"ec"),
  1437 => (x"87",x"c5",x"d5",x"49"),
  1438 => (x"ff",x"1e",x"4f",x"26"),
  1439 => (x"ff",x"c3",x"4a",x"d4"),
  1440 => (x"48",x"d0",x"ff",x"7a"),
  1441 => (x"de",x"78",x"e1",x"c0"),
  1442 => (x"48",x"7a",x"71",x"7a"),
  1443 => (x"70",x"28",x"b7",x"c8"),
  1444 => (x"d0",x"48",x"71",x"7a"),
  1445 => (x"7a",x"70",x"28",x"b7"),
  1446 => (x"b7",x"d8",x"48",x"71"),
  1447 => (x"ff",x"7a",x"70",x"28"),
  1448 => (x"e0",x"c0",x"48",x"d0"),
  1449 => (x"0e",x"4f",x"26",x"78"),
  1450 => (x"5d",x"5c",x"5b",x"5e"),
  1451 => (x"71",x"86",x"f4",x"0e"),
  1452 => (x"91",x"cc",x"49",x"4d"),
  1453 => (x"81",x"f8",x"f1",x"c1"),
  1454 => (x"ca",x"4a",x"a1",x"c8"),
  1455 => (x"a6",x"c4",x"7e",x"a1"),
  1456 => (x"d4",x"f5",x"c2",x"48"),
  1457 => (x"97",x"6e",x"78",x"bf"),
  1458 => (x"66",x"c4",x"4b",x"bf"),
  1459 => (x"12",x"2c",x"73",x"4c"),
  1460 => (x"58",x"a6",x"cc",x"48"),
  1461 => (x"84",x"c1",x"9c",x"70"),
  1462 => (x"69",x"97",x"81",x"c9"),
  1463 => (x"04",x"ac",x"b7",x"49"),
  1464 => (x"4c",x"c0",x"87",x"c2"),
  1465 => (x"4a",x"bf",x"97",x"6e"),
  1466 => (x"72",x"49",x"66",x"c8"),
  1467 => (x"c4",x"b9",x"ff",x"31"),
  1468 => (x"48",x"74",x"99",x"66"),
  1469 => (x"4a",x"70",x"30",x"72"),
  1470 => (x"d8",x"f5",x"c2",x"b1"),
  1471 => (x"f9",x"fd",x"71",x"59"),
  1472 => (x"c2",x"1e",x"c7",x"87"),
  1473 => (x"1e",x"bf",x"e8",x"f6"),
  1474 => (x"1e",x"f8",x"f1",x"c1"),
  1475 => (x"97",x"d8",x"f5",x"c2"),
  1476 => (x"f4",x"c1",x"49",x"bf"),
  1477 => (x"c0",x"49",x"75",x"87"),
  1478 => (x"e8",x"87",x"e1",x"f3"),
  1479 => (x"26",x"4d",x"26",x"8e"),
  1480 => (x"26",x"4b",x"26",x"4c"),
  1481 => (x"1e",x"73",x"1e",x"4f"),
  1482 => (x"fd",x"49",x"4b",x"71"),
  1483 => (x"49",x"73",x"87",x"f9"),
  1484 => (x"26",x"87",x"f4",x"fd"),
  1485 => (x"1e",x"4f",x"26",x"4b"),
  1486 => (x"4b",x"71",x"1e",x"73"),
  1487 => (x"02",x"4a",x"a3",x"c2"),
  1488 => (x"8a",x"c1",x"87",x"d6"),
  1489 => (x"87",x"e2",x"c0",x"05"),
  1490 => (x"bf",x"e8",x"f6",x"c2"),
  1491 => (x"48",x"87",x"db",x"02"),
  1492 => (x"f6",x"c2",x"88",x"c1"),
  1493 => (x"87",x"d2",x"58",x"ec"),
  1494 => (x"bf",x"ec",x"f6",x"c2"),
  1495 => (x"c2",x"87",x"cb",x"02"),
  1496 => (x"48",x"bf",x"e8",x"f6"),
  1497 => (x"f6",x"c2",x"80",x"c1"),
  1498 => (x"1e",x"c7",x"58",x"ec"),
  1499 => (x"bf",x"e8",x"f6",x"c2"),
  1500 => (x"f8",x"f1",x"c1",x"1e"),
  1501 => (x"d8",x"f5",x"c2",x"1e"),
  1502 => (x"cc",x"49",x"bf",x"97"),
  1503 => (x"c0",x"49",x"73",x"87"),
  1504 => (x"f4",x"87",x"f9",x"f1"),
  1505 => (x"26",x"4b",x"26",x"8e"),
  1506 => (x"5b",x"5e",x"0e",x"4f"),
  1507 => (x"ff",x"0e",x"5d",x"5c"),
  1508 => (x"e8",x"c0",x"86",x"cc"),
  1509 => (x"a6",x"cc",x"59",x"a6"),
  1510 => (x"c4",x"78",x"c0",x"48"),
  1511 => (x"c4",x"78",x"c0",x"80"),
  1512 => (x"c4",x"78",x"c0",x"80"),
  1513 => (x"66",x"c8",x"c1",x"80"),
  1514 => (x"c1",x"80",x"c4",x"78"),
  1515 => (x"c1",x"80",x"c4",x"78"),
  1516 => (x"ec",x"f6",x"c2",x"78"),
  1517 => (x"ff",x"78",x"c1",x"48"),
  1518 => (x"ff",x"87",x"e4",x"df"),
  1519 => (x"ff",x"87",x"fd",x"df"),
  1520 => (x"70",x"87",x"d1",x"df"),
  1521 => (x"ad",x"fb",x"c0",x"4d"),
  1522 => (x"87",x"f3",x"c1",x"02"),
  1523 => (x"05",x"66",x"e4",x"c0"),
  1524 => (x"c1",x"87",x"e8",x"c1"),
  1525 => (x"c4",x"4a",x"66",x"c4"),
  1526 => (x"c1",x"7e",x"6a",x"82"),
  1527 => (x"6e",x"48",x"e0",x"ca"),
  1528 => (x"20",x"41",x"20",x"49"),
  1529 => (x"c1",x"51",x"10",x"41"),
  1530 => (x"c1",x"48",x"66",x"c4"),
  1531 => (x"6a",x"78",x"e1",x"d8"),
  1532 => (x"75",x"81",x"c7",x"49"),
  1533 => (x"66",x"c4",x"c1",x"51"),
  1534 => (x"c1",x"81",x"c8",x"49"),
  1535 => (x"48",x"a6",x"dc",x"51"),
  1536 => (x"c4",x"c1",x"78",x"c2"),
  1537 => (x"81",x"c9",x"49",x"66"),
  1538 => (x"c4",x"c1",x"51",x"c0"),
  1539 => (x"81",x"ca",x"49",x"66"),
  1540 => (x"1e",x"c1",x"51",x"c0"),
  1541 => (x"49",x"6a",x"1e",x"d8"),
  1542 => (x"de",x"ff",x"81",x"c8"),
  1543 => (x"86",x"c8",x"87",x"f2"),
  1544 => (x"48",x"66",x"c8",x"c1"),
  1545 => (x"c7",x"01",x"a8",x"c0"),
  1546 => (x"48",x"a6",x"d4",x"87"),
  1547 => (x"87",x"cf",x"78",x"c1"),
  1548 => (x"48",x"66",x"c8",x"c1"),
  1549 => (x"a6",x"dc",x"88",x"c1"),
  1550 => (x"ff",x"87",x"c4",x"58"),
  1551 => (x"75",x"87",x"fd",x"dd"),
  1552 => (x"f2",x"cb",x"02",x"9d"),
  1553 => (x"48",x"66",x"d4",x"87"),
  1554 => (x"a8",x"66",x"cc",x"c1"),
  1555 => (x"87",x"e7",x"cb",x"03"),
  1556 => (x"dc",x"ff",x"7e",x"c0"),
  1557 => (x"4d",x"70",x"87",x"fe"),
  1558 => (x"88",x"c6",x"c1",x"48"),
  1559 => (x"70",x"58",x"a6",x"c8"),
  1560 => (x"d6",x"c1",x"02",x"98"),
  1561 => (x"88",x"c9",x"48",x"87"),
  1562 => (x"70",x"58",x"a6",x"c8"),
  1563 => (x"d8",x"c5",x"02",x"98"),
  1564 => (x"88",x"c1",x"48",x"87"),
  1565 => (x"70",x"58",x"a6",x"c8"),
  1566 => (x"f8",x"c2",x"02",x"98"),
  1567 => (x"88",x"c3",x"48",x"87"),
  1568 => (x"70",x"58",x"a6",x"c8"),
  1569 => (x"87",x"cf",x"02",x"98"),
  1570 => (x"c8",x"88",x"c1",x"48"),
  1571 => (x"98",x"70",x"58",x"a6"),
  1572 => (x"87",x"f5",x"c4",x"02"),
  1573 => (x"c0",x"87",x"ff",x"c9"),
  1574 => (x"db",x"ff",x"7e",x"f0"),
  1575 => (x"4d",x"70",x"87",x"f6"),
  1576 => (x"02",x"ad",x"ec",x"c0"),
  1577 => (x"7e",x"75",x"87",x"c2"),
  1578 => (x"02",x"ad",x"ec",x"c0"),
  1579 => (x"db",x"ff",x"87",x"cd"),
  1580 => (x"4d",x"70",x"87",x"e2"),
  1581 => (x"05",x"ad",x"ec",x"c0"),
  1582 => (x"c0",x"87",x"f3",x"ff"),
  1583 => (x"c1",x"05",x"66",x"e4"),
  1584 => (x"ec",x"c0",x"87",x"ea"),
  1585 => (x"87",x"c4",x"02",x"ad"),
  1586 => (x"87",x"c8",x"db",x"ff"),
  1587 => (x"1e",x"ca",x"1e",x"c0"),
  1588 => (x"cc",x"4b",x"66",x"dc"),
  1589 => (x"66",x"cc",x"c1",x"93"),
  1590 => (x"4c",x"a3",x"c4",x"83"),
  1591 => (x"db",x"ff",x"49",x"6c"),
  1592 => (x"1e",x"c1",x"87",x"ee"),
  1593 => (x"49",x"6c",x"1e",x"de"),
  1594 => (x"87",x"e4",x"db",x"ff"),
  1595 => (x"d8",x"c1",x"86",x"d0"),
  1596 => (x"a3",x"c8",x"7b",x"e1"),
  1597 => (x"51",x"66",x"dc",x"49"),
  1598 => (x"c0",x"49",x"a3",x"c9"),
  1599 => (x"ca",x"51",x"66",x"e0"),
  1600 => (x"51",x"6e",x"49",x"a3"),
  1601 => (x"c1",x"48",x"66",x"dc"),
  1602 => (x"a6",x"e0",x"c0",x"80"),
  1603 => (x"48",x"66",x"d4",x"58"),
  1604 => (x"04",x"a8",x"66",x"d8"),
  1605 => (x"66",x"d4",x"87",x"cb"),
  1606 => (x"d8",x"80",x"c1",x"48"),
  1607 => (x"fb",x"c7",x"58",x"a6"),
  1608 => (x"48",x"66",x"d8",x"87"),
  1609 => (x"a6",x"dc",x"88",x"c1"),
  1610 => (x"87",x"f0",x"c7",x"58"),
  1611 => (x"87",x"cc",x"da",x"ff"),
  1612 => (x"e7",x"c7",x"4d",x"70"),
  1613 => (x"c2",x"dc",x"ff",x"87"),
  1614 => (x"58",x"a6",x"d0",x"87"),
  1615 => (x"06",x"a8",x"66",x"d0"),
  1616 => (x"d0",x"87",x"c6",x"c0"),
  1617 => (x"66",x"cc",x"48",x"a6"),
  1618 => (x"ee",x"db",x"ff",x"78"),
  1619 => (x"a8",x"ec",x"c0",x"87"),
  1620 => (x"87",x"f5",x"c1",x"05"),
  1621 => (x"05",x"66",x"e4",x"c0"),
  1622 => (x"d4",x"87",x"e5",x"c1"),
  1623 => (x"91",x"cc",x"49",x"66"),
  1624 => (x"81",x"66",x"c4",x"c1"),
  1625 => (x"6a",x"4a",x"a1",x"c4"),
  1626 => (x"4a",x"a1",x"c8",x"4c"),
  1627 => (x"c1",x"52",x"66",x"cc"),
  1628 => (x"ff",x"79",x"d9",x"d9"),
  1629 => (x"70",x"87",x"dd",x"d8"),
  1630 => (x"da",x"02",x"9d",x"4d"),
  1631 => (x"ad",x"fb",x"c0",x"87"),
  1632 => (x"75",x"87",x"d4",x"02"),
  1633 => (x"cb",x"d8",x"ff",x"54"),
  1634 => (x"9d",x"4d",x"70",x"87"),
  1635 => (x"87",x"c7",x"c0",x"02"),
  1636 => (x"05",x"ad",x"fb",x"c0"),
  1637 => (x"c0",x"87",x"ec",x"ff"),
  1638 => (x"c1",x"c2",x"54",x"e0"),
  1639 => (x"7c",x"97",x"c0",x"54"),
  1640 => (x"d8",x"48",x"66",x"d4"),
  1641 => (x"c0",x"04",x"a8",x"66"),
  1642 => (x"66",x"d4",x"87",x"cb"),
  1643 => (x"d8",x"80",x"c1",x"48"),
  1644 => (x"e7",x"c5",x"58",x"a6"),
  1645 => (x"48",x"66",x"d8",x"87"),
  1646 => (x"a6",x"dc",x"88",x"c1"),
  1647 => (x"87",x"dc",x"c5",x"58"),
  1648 => (x"87",x"f8",x"d7",x"ff"),
  1649 => (x"d3",x"c5",x"4d",x"70"),
  1650 => (x"48",x"66",x"cc",x"87"),
  1651 => (x"a8",x"66",x"e4",x"c0"),
  1652 => (x"87",x"f4",x"c4",x"05"),
  1653 => (x"48",x"a6",x"e8",x"c0"),
  1654 => (x"d9",x"ff",x"78",x"c0"),
  1655 => (x"7e",x"70",x"87",x"dd"),
  1656 => (x"87",x"d7",x"d9",x"ff"),
  1657 => (x"58",x"a6",x"f0",x"c0"),
  1658 => (x"05",x"a8",x"ec",x"c0"),
  1659 => (x"a6",x"87",x"c7",x"c0"),
  1660 => (x"c0",x"78",x"6e",x"48"),
  1661 => (x"d6",x"ff",x"87",x"c4"),
  1662 => (x"66",x"d4",x"87",x"da"),
  1663 => (x"c1",x"91",x"cc",x"49"),
  1664 => (x"71",x"48",x"66",x"c4"),
  1665 => (x"58",x"a6",x"c8",x"80"),
  1666 => (x"c8",x"4a",x"66",x"c4"),
  1667 => (x"49",x"66",x"c4",x"82"),
  1668 => (x"51",x"6e",x"81",x"ca"),
  1669 => (x"49",x"66",x"ec",x"c0"),
  1670 => (x"89",x"6e",x"81",x"c1"),
  1671 => (x"30",x"71",x"48",x"c1"),
  1672 => (x"89",x"c1",x"49",x"70"),
  1673 => (x"c2",x"7a",x"97",x"71"),
  1674 => (x"49",x"bf",x"d4",x"f5"),
  1675 => (x"6a",x"97",x"29",x"6e"),
  1676 => (x"98",x"71",x"48",x"4a"),
  1677 => (x"58",x"a6",x"f4",x"c0"),
  1678 => (x"c4",x"48",x"66",x"c4"),
  1679 => (x"58",x"a6",x"cc",x"80"),
  1680 => (x"4c",x"bf",x"66",x"c8"),
  1681 => (x"48",x"66",x"e4",x"c0"),
  1682 => (x"02",x"a8",x"66",x"cc"),
  1683 => (x"c0",x"87",x"c5",x"c0"),
  1684 => (x"87",x"c2",x"c0",x"7e"),
  1685 => (x"1e",x"6e",x"7e",x"c1"),
  1686 => (x"74",x"1e",x"e0",x"c0"),
  1687 => (x"ef",x"d5",x"ff",x"49"),
  1688 => (x"70",x"86",x"c8",x"87"),
  1689 => (x"ad",x"b7",x"c0",x"4d"),
  1690 => (x"87",x"d4",x"c1",x"06"),
  1691 => (x"66",x"c8",x"84",x"75"),
  1692 => (x"e0",x"c0",x"49",x"bf"),
  1693 => (x"4b",x"89",x"74",x"81"),
  1694 => (x"4a",x"ec",x"ca",x"c1"),
  1695 => (x"e1",x"de",x"fe",x"71"),
  1696 => (x"74",x"84",x"c2",x"87"),
  1697 => (x"66",x"e8",x"c0",x"7e"),
  1698 => (x"c0",x"80",x"c1",x"48"),
  1699 => (x"c0",x"58",x"a6",x"ec"),
  1700 => (x"c1",x"49",x"66",x"f0"),
  1701 => (x"02",x"a9",x"70",x"81"),
  1702 => (x"c0",x"87",x"c5",x"c0"),
  1703 => (x"87",x"c2",x"c0",x"4c"),
  1704 => (x"1e",x"74",x"4c",x"c1"),
  1705 => (x"49",x"bf",x"66",x"cc"),
  1706 => (x"c4",x"81",x"e0",x"c0"),
  1707 => (x"1e",x"71",x"89",x"66"),
  1708 => (x"ff",x"49",x"66",x"c8"),
  1709 => (x"c8",x"87",x"d9",x"d4"),
  1710 => (x"a8",x"b7",x"c0",x"86"),
  1711 => (x"87",x"c5",x"ff",x"01"),
  1712 => (x"02",x"66",x"e8",x"c0"),
  1713 => (x"c4",x"87",x"d3",x"c0"),
  1714 => (x"81",x"c9",x"49",x"66"),
  1715 => (x"51",x"66",x"e8",x"c0"),
  1716 => (x"c1",x"48",x"66",x"c4"),
  1717 => (x"c0",x"78",x"e7",x"da"),
  1718 => (x"66",x"c4",x"87",x"ce"),
  1719 => (x"c2",x"81",x"c9",x"49"),
  1720 => (x"48",x"66",x"c4",x"51"),
  1721 => (x"78",x"e5",x"dc",x"c1"),
  1722 => (x"d8",x"48",x"66",x"d4"),
  1723 => (x"c0",x"04",x"a8",x"66"),
  1724 => (x"66",x"d4",x"87",x"cb"),
  1725 => (x"d8",x"80",x"c1",x"48"),
  1726 => (x"d1",x"c0",x"58",x"a6"),
  1727 => (x"48",x"66",x"d8",x"87"),
  1728 => (x"a6",x"dc",x"88",x"c1"),
  1729 => (x"87",x"c6",x"c0",x"58"),
  1730 => (x"87",x"f0",x"d2",x"ff"),
  1731 => (x"a6",x"cc",x"4d",x"70"),
  1732 => (x"c0",x"78",x"c0",x"48"),
  1733 => (x"d2",x"ff",x"87",x"c6"),
  1734 => (x"4d",x"70",x"87",x"e2"),
  1735 => (x"48",x"66",x"e0",x"c0"),
  1736 => (x"e4",x"c0",x"80",x"c1"),
  1737 => (x"9d",x"75",x"58",x"a6"),
  1738 => (x"87",x"cb",x"c0",x"02"),
  1739 => (x"c1",x"48",x"66",x"d4"),
  1740 => (x"04",x"a8",x"66",x"cc"),
  1741 => (x"d4",x"87",x"d9",x"f4"),
  1742 => (x"a8",x"c7",x"48",x"66"),
  1743 => (x"87",x"e1",x"c0",x"03"),
  1744 => (x"c2",x"4c",x"66",x"d4"),
  1745 => (x"c0",x"48",x"ec",x"f6"),
  1746 => (x"cc",x"49",x"74",x"78"),
  1747 => (x"66",x"c4",x"c1",x"91"),
  1748 => (x"4a",x"a1",x"c4",x"81"),
  1749 => (x"52",x"c0",x"4a",x"6a"),
  1750 => (x"c7",x"84",x"c1",x"79"),
  1751 => (x"e2",x"ff",x"04",x"ac"),
  1752 => (x"66",x"e4",x"c0",x"87"),
  1753 => (x"87",x"e2",x"c0",x"02"),
  1754 => (x"49",x"66",x"c4",x"c1"),
  1755 => (x"c1",x"81",x"d4",x"c1"),
  1756 => (x"c1",x"4a",x"66",x"c4"),
  1757 => (x"52",x"c0",x"82",x"dc"),
  1758 => (x"79",x"d9",x"d9",x"c1"),
  1759 => (x"49",x"66",x"c4",x"c1"),
  1760 => (x"c1",x"81",x"d8",x"c1"),
  1761 => (x"c0",x"79",x"f0",x"ca"),
  1762 => (x"c4",x"c1",x"87",x"d6"),
  1763 => (x"d4",x"c1",x"49",x"66"),
  1764 => (x"66",x"c4",x"c1",x"81"),
  1765 => (x"82",x"d8",x"c1",x"4a"),
  1766 => (x"7a",x"f8",x"ca",x"c1"),
  1767 => (x"79",x"d0",x"d9",x"c1"),
  1768 => (x"49",x"66",x"c4",x"c1"),
  1769 => (x"c1",x"81",x"e0",x"c1"),
  1770 => (x"ff",x"79",x"f7",x"dc"),
  1771 => (x"d0",x"87",x"c4",x"d0"),
  1772 => (x"cc",x"ff",x"48",x"66"),
  1773 => (x"26",x"4d",x"26",x"8e"),
  1774 => (x"26",x"4b",x"26",x"4c"),
  1775 => (x"1e",x"c7",x"1e",x"4f"),
  1776 => (x"bf",x"e8",x"f6",x"c2"),
  1777 => (x"f8",x"f1",x"c1",x"1e"),
  1778 => (x"d8",x"f5",x"c2",x"1e"),
  1779 => (x"ee",x"49",x"bf",x"97"),
  1780 => (x"f1",x"c1",x"87",x"f7"),
  1781 => (x"e1",x"c0",x"49",x"f8"),
  1782 => (x"8e",x"f4",x"87",x"f0"),
  1783 => (x"c1",x"1e",x"4f",x"26"),
  1784 => (x"c0",x"48",x"ec",x"f1"),
  1785 => (x"e4",x"f3",x"c1",x"50"),
  1786 => (x"d4",x"ff",x"49",x"bf"),
  1787 => (x"48",x"c0",x"87",x"fc"),
  1788 => (x"73",x"1e",x"4f",x"26"),
  1789 => (x"87",x"ce",x"c7",x"1e"),
  1790 => (x"48",x"f4",x"f6",x"c2"),
  1791 => (x"d4",x"ff",x"50",x"c0"),
  1792 => (x"78",x"ff",x"c3",x"48"),
  1793 => (x"49",x"c0",x"cb",x"c1"),
  1794 => (x"87",x"fd",x"d6",x"fe"),
  1795 => (x"87",x"d0",x"e2",x"fe"),
  1796 => (x"cd",x"02",x"98",x"70"),
  1797 => (x"ee",x"eb",x"fe",x"87"),
  1798 => (x"02",x"98",x"70",x"87"),
  1799 => (x"4a",x"c1",x"87",x"c4"),
  1800 => (x"4a",x"c0",x"87",x"c2"),
  1801 => (x"c8",x"02",x"9a",x"72"),
  1802 => (x"cc",x"cb",x"c1",x"87"),
  1803 => (x"d8",x"d6",x"fe",x"49"),
  1804 => (x"e8",x"f6",x"c2",x"87"),
  1805 => (x"c2",x"78",x"c0",x"48"),
  1806 => (x"c0",x"48",x"d8",x"f5"),
  1807 => (x"fc",x"fd",x"49",x"50"),
  1808 => (x"87",x"da",x"fe",x"87"),
  1809 => (x"02",x"9b",x"4b",x"70"),
  1810 => (x"f3",x"c1",x"87",x"cf"),
  1811 => (x"49",x"c7",x"5b",x"d4"),
  1812 => (x"c1",x"87",x"e9",x"de"),
  1813 => (x"c4",x"e0",x"c0",x"49"),
  1814 => (x"87",x"f3",x"c2",x"87"),
  1815 => (x"87",x"ca",x"e1",x"c0"),
  1816 => (x"87",x"dc",x"ef",x"c0"),
  1817 => (x"26",x"87",x"f5",x"ff"),
  1818 => (x"00",x"4f",x"26",x"4b"),
  1819 => (x"00",x"00",x"00",x"00"),
  1820 => (x"00",x"00",x"00",x"00"),
  1821 => (x"00",x"00",x"00",x"01"),
  1822 => (x"00",x"00",x"13",x"65"),
  1823 => (x"00",x"00",x"2d",x"c0"),
  1824 => (x"94",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"13",x"65"),
  1826 => (x"00",x"00",x"2d",x"de"),
  1827 => (x"94",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"13",x"65"),
  1829 => (x"00",x"00",x"2d",x"fc"),
  1830 => (x"94",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"13",x"65"),
  1832 => (x"00",x"00",x"2e",x"1a"),
  1833 => (x"94",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"13",x"65"),
  1835 => (x"00",x"00",x"2e",x"38"),
  1836 => (x"94",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"13",x"65"),
  1838 => (x"00",x"00",x"2e",x"56"),
  1839 => (x"94",x"00",x"00",x"00"),
  1840 => (x"00",x"00",x"13",x"65"),
  1841 => (x"00",x"00",x"2e",x"74"),
  1842 => (x"94",x"00",x"00",x"00"),
  1843 => (x"00",x"00",x"16",x"59"),
  1844 => (x"00",x"00",x"00",x"00"),
  1845 => (x"94",x"00",x"00",x"00"),
  1846 => (x"00",x"00",x"14",x"0b"),
  1847 => (x"00",x"00",x"00",x"00"),
  1848 => (x"94",x"00",x"00",x"00"),
  1849 => (x"00",x"00",x"12",x"d0"),
  1850 => (x"db",x"86",x"fc",x"1e"),
  1851 => (x"fc",x"7e",x"70",x"87"),
  1852 => (x"1e",x"4f",x"26",x"8e"),
  1853 => (x"c0",x"48",x"f0",x"fe"),
  1854 => (x"79",x"09",x"cd",x"78"),
  1855 => (x"1e",x"4f",x"26",x"09"),
  1856 => (x"49",x"e8",x"f3",x"c1"),
  1857 => (x"4f",x"26",x"87",x"ed"),
  1858 => (x"bf",x"f0",x"fe",x"1e"),
  1859 => (x"1e",x"4f",x"26",x"48"),
  1860 => (x"c1",x"48",x"f0",x"fe"),
  1861 => (x"1e",x"4f",x"26",x"78"),
  1862 => (x"c0",x"48",x"f0",x"fe"),
  1863 => (x"1e",x"4f",x"26",x"78"),
  1864 => (x"52",x"c0",x"4a",x"71"),
  1865 => (x"0e",x"4f",x"26",x"51"),
  1866 => (x"5d",x"5c",x"5b",x"5e"),
  1867 => (x"71",x"86",x"f4",x"0e"),
  1868 => (x"7e",x"6d",x"97",x"4d"),
  1869 => (x"97",x"4c",x"a5",x"c1"),
  1870 => (x"a6",x"c8",x"48",x"6c"),
  1871 => (x"c4",x"48",x"6e",x"58"),
  1872 => (x"c5",x"05",x"a8",x"66"),
  1873 => (x"c0",x"48",x"ff",x"87"),
  1874 => (x"ca",x"ff",x"87",x"e6"),
  1875 => (x"49",x"a5",x"c2",x"87"),
  1876 => (x"71",x"4b",x"6c",x"97"),
  1877 => (x"6b",x"97",x"4b",x"a3"),
  1878 => (x"7e",x"6c",x"97",x"4b"),
  1879 => (x"80",x"c1",x"48",x"6e"),
  1880 => (x"c7",x"58",x"a6",x"c8"),
  1881 => (x"58",x"a6",x"cc",x"98"),
  1882 => (x"fe",x"7c",x"97",x"70"),
  1883 => (x"48",x"73",x"87",x"e1"),
  1884 => (x"4d",x"26",x"8e",x"f4"),
  1885 => (x"4b",x"26",x"4c",x"26"),
  1886 => (x"73",x"1e",x"4f",x"26"),
  1887 => (x"fe",x"86",x"f4",x"1e"),
  1888 => (x"bf",x"e0",x"87",x"d5"),
  1889 => (x"e0",x"c0",x"49",x"4b"),
  1890 => (x"c0",x"02",x"99",x"c0"),
  1891 => (x"4a",x"73",x"87",x"ea"),
  1892 => (x"c2",x"9a",x"ff",x"c3"),
  1893 => (x"bf",x"97",x"e8",x"fa"),
  1894 => (x"ea",x"fa",x"c2",x"49"),
  1895 => (x"c2",x"51",x"72",x"81"),
  1896 => (x"bf",x"97",x"e8",x"fa"),
  1897 => (x"c1",x"48",x"6e",x"7e"),
  1898 => (x"58",x"a6",x"c8",x"80"),
  1899 => (x"a6",x"cc",x"98",x"c7"),
  1900 => (x"e8",x"fa",x"c2",x"58"),
  1901 => (x"50",x"66",x"c8",x"48"),
  1902 => (x"70",x"87",x"cd",x"fd"),
  1903 => (x"87",x"cf",x"fd",x"7e"),
  1904 => (x"4b",x"26",x"8e",x"f4"),
  1905 => (x"c2",x"1e",x"4f",x"26"),
  1906 => (x"fd",x"49",x"e8",x"fa"),
  1907 => (x"f5",x"c1",x"87",x"d1"),
  1908 => (x"de",x"fc",x"49",x"fa"),
  1909 => (x"87",x"e8",x"c4",x"87"),
  1910 => (x"5e",x"0e",x"4f",x"26"),
  1911 => (x"0e",x"5d",x"5c",x"5b"),
  1912 => (x"7e",x"71",x"86",x"fc"),
  1913 => (x"c2",x"4d",x"d4",x"ff"),
  1914 => (x"fc",x"49",x"e8",x"fa"),
  1915 => (x"4b",x"70",x"87",x"f9"),
  1916 => (x"04",x"ab",x"b7",x"c0"),
  1917 => (x"c3",x"87",x"f5",x"c2"),
  1918 => (x"c9",x"05",x"ab",x"f0"),
  1919 => (x"f8",x"fa",x"c1",x"87"),
  1920 => (x"c2",x"78",x"c1",x"48"),
  1921 => (x"e0",x"c3",x"87",x"d6"),
  1922 => (x"87",x"c9",x"05",x"ab"),
  1923 => (x"48",x"fc",x"fa",x"c1"),
  1924 => (x"c7",x"c2",x"78",x"c1"),
  1925 => (x"fc",x"fa",x"c1",x"87"),
  1926 => (x"87",x"c6",x"02",x"bf"),
  1927 => (x"4c",x"a3",x"c0",x"c2"),
  1928 => (x"4c",x"73",x"87",x"c2"),
  1929 => (x"bf",x"f8",x"fa",x"c1"),
  1930 => (x"87",x"e0",x"c0",x"02"),
  1931 => (x"b7",x"c4",x"49",x"74"),
  1932 => (x"fb",x"c1",x"91",x"29"),
  1933 => (x"4a",x"74",x"81",x"c0"),
  1934 => (x"92",x"c2",x"9a",x"cf"),
  1935 => (x"30",x"72",x"48",x"c1"),
  1936 => (x"ba",x"ff",x"4a",x"70"),
  1937 => (x"98",x"69",x"48",x"72"),
  1938 => (x"87",x"db",x"79",x"70"),
  1939 => (x"b7",x"c4",x"49",x"74"),
  1940 => (x"fb",x"c1",x"91",x"29"),
  1941 => (x"4a",x"74",x"81",x"c0"),
  1942 => (x"92",x"c2",x"9a",x"cf"),
  1943 => (x"30",x"72",x"48",x"c3"),
  1944 => (x"69",x"48",x"4a",x"70"),
  1945 => (x"6e",x"79",x"70",x"b0"),
  1946 => (x"87",x"e4",x"c0",x"05"),
  1947 => (x"c8",x"48",x"d0",x"ff"),
  1948 => (x"7d",x"c5",x"78",x"e1"),
  1949 => (x"bf",x"fc",x"fa",x"c1"),
  1950 => (x"c3",x"87",x"c3",x"02"),
  1951 => (x"fa",x"c1",x"7d",x"e0"),
  1952 => (x"c3",x"02",x"bf",x"f8"),
  1953 => (x"7d",x"f0",x"c3",x"87"),
  1954 => (x"d0",x"ff",x"7d",x"73"),
  1955 => (x"78",x"e0",x"c0",x"48"),
  1956 => (x"48",x"fc",x"fa",x"c1"),
  1957 => (x"fa",x"c1",x"78",x"c0"),
  1958 => (x"78",x"c0",x"48",x"f8"),
  1959 => (x"49",x"e8",x"fa",x"c2"),
  1960 => (x"70",x"87",x"c4",x"fa"),
  1961 => (x"ab",x"b7",x"c0",x"4b"),
  1962 => (x"87",x"cb",x"fd",x"03"),
  1963 => (x"8e",x"fc",x"48",x"c0"),
  1964 => (x"4c",x"26",x"4d",x"26"),
  1965 => (x"4f",x"26",x"4b",x"26"),
  1966 => (x"00",x"00",x"00",x"00"),
  1967 => (x"00",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"84",x"84",x"84",x"84"),
  1970 => (x"84",x"84",x"84",x"84"),
  1971 => (x"84",x"84",x"84",x"84"),
  1972 => (x"84",x"84",x"84",x"84"),
  1973 => (x"84",x"84",x"84",x"84"),
  1974 => (x"84",x"84",x"84",x"84"),
  1975 => (x"84",x"84",x"84",x"84"),
  1976 => (x"84",x"84",x"84",x"84"),
  1977 => (x"84",x"84",x"84",x"84"),
  1978 => (x"84",x"84",x"84",x"84"),
  1979 => (x"84",x"84",x"84",x"84"),
  1980 => (x"84",x"84",x"84",x"84"),
  1981 => (x"84",x"84",x"84",x"84"),
  1982 => (x"84",x"84",x"84",x"84"),
  1983 => (x"84",x"84",x"84",x"84"),
  1984 => (x"72",x"4a",x"c0",x"1e"),
  1985 => (x"c1",x"91",x"c4",x"49"),
  1986 => (x"c0",x"81",x"c0",x"fb"),
  1987 => (x"d0",x"82",x"c1",x"79"),
  1988 => (x"ee",x"04",x"aa",x"b7"),
  1989 => (x"0e",x"4f",x"26",x"87"),
  1990 => (x"5d",x"5c",x"5b",x"5e"),
  1991 => (x"f7",x"4d",x"71",x"0e"),
  1992 => (x"4a",x"75",x"87",x"f5"),
  1993 => (x"92",x"2a",x"b7",x"c4"),
  1994 => (x"82",x"c0",x"fb",x"c1"),
  1995 => (x"9c",x"cf",x"4c",x"75"),
  1996 => (x"49",x"6a",x"94",x"c2"),
  1997 => (x"c3",x"2b",x"74",x"4b"),
  1998 => (x"74",x"48",x"c2",x"9b"),
  1999 => (x"ff",x"4c",x"70",x"30"),
  2000 => (x"71",x"48",x"74",x"bc"),
  2001 => (x"f7",x"7a",x"70",x"98"),
  2002 => (x"48",x"73",x"87",x"c5"),
  2003 => (x"4c",x"26",x"4d",x"26"),
  2004 => (x"4f",x"26",x"4b",x"26"),
  2005 => (x"48",x"d0",x"ff",x"1e"),
  2006 => (x"71",x"78",x"e1",x"c8"),
  2007 => (x"08",x"d4",x"ff",x"48"),
  2008 => (x"1e",x"4f",x"26",x"78"),
  2009 => (x"c8",x"48",x"d0",x"ff"),
  2010 => (x"48",x"71",x"78",x"e1"),
  2011 => (x"78",x"08",x"d4",x"ff"),
  2012 => (x"ff",x"48",x"66",x"c4"),
  2013 => (x"26",x"78",x"08",x"d4"),
  2014 => (x"4a",x"71",x"1e",x"4f"),
  2015 => (x"1e",x"49",x"66",x"c4"),
  2016 => (x"de",x"ff",x"49",x"72"),
  2017 => (x"48",x"d0",x"ff",x"87"),
  2018 => (x"fc",x"78",x"e0",x"c0"),
  2019 => (x"1e",x"4f",x"26",x"8e"),
  2020 => (x"4b",x"71",x"1e",x"73"),
  2021 => (x"1e",x"49",x"66",x"c8"),
  2022 => (x"e0",x"c1",x"4a",x"73"),
  2023 => (x"d8",x"ff",x"49",x"a2"),
  2024 => (x"26",x"8e",x"fc",x"87"),
  2025 => (x"1e",x"4f",x"26",x"4b"),
  2026 => (x"c8",x"48",x"d0",x"ff"),
  2027 => (x"48",x"71",x"78",x"c9"),
  2028 => (x"78",x"08",x"d4",x"ff"),
  2029 => (x"71",x"1e",x"4f",x"26"),
  2030 => (x"87",x"eb",x"49",x"4a"),
  2031 => (x"c8",x"48",x"d0",x"ff"),
  2032 => (x"1e",x"4f",x"26",x"78"),
  2033 => (x"4b",x"71",x"1e",x"73"),
  2034 => (x"bf",x"c0",x"fb",x"c2"),
  2035 => (x"c2",x"87",x"c3",x"02"),
  2036 => (x"d0",x"ff",x"87",x"eb"),
  2037 => (x"78",x"c9",x"c8",x"48"),
  2038 => (x"e0",x"c0",x"48",x"73"),
  2039 => (x"08",x"d4",x"ff",x"b0"),
  2040 => (x"f4",x"fa",x"c2",x"78"),
  2041 => (x"c8",x"78",x"c0",x"48"),
  2042 => (x"87",x"c5",x"02",x"66"),
  2043 => (x"c2",x"49",x"ff",x"c3"),
  2044 => (x"c2",x"49",x"c0",x"87"),
  2045 => (x"cc",x"59",x"fc",x"fa"),
  2046 => (x"87",x"c6",x"02",x"66"),
  2047 => (x"4a",x"d5",x"d5",x"c5"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

