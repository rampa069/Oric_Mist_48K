library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ecc0c387",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49ecc0c3",
    18 => x"48c4e8c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"c3e8c287",
    25 => x"ffe7c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"eec187f7",
    29 => x"e8c287d1",
    30 => x"e8c24dc3",
    31 => x"ad744cc3",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"5c5b5e0e",
    36 => x"86f00e5d",
    37 => x"a6c44cc0",
    38 => x"c078c048",
    39 => x"c04ba6e4",
    40 => x"484966e0",
    41 => x"e4c080c1",
    42 => x"481158a6",
    43 => x"7058a6c4",
    44 => x"f6c30298",
    45 => x"0266c487",
    46 => x"c487c6c3",
    47 => x"78c048a6",
    48 => x"f0c04a6e",
    49 => x"dac2028a",
    50 => x"8af3c087",
    51 => x"87dbc202",
    52 => x"dc028ac1",
    53 => x"028ac887",
    54 => x"c487c8c2",
    55 => x"87d1028a",
    56 => x"c1028ac3",
    57 => x"8ac287eb",
    58 => x"c387c602",
    59 => x"c9c2058a",
    60 => x"7383c487",
    61 => x"6989c449",
    62 => x"c1026e7e",
    63 => x"a6c887c8",
    64 => x"c478c048",
    65 => x"cc78c080",
    66 => x"4a6e4d66",
    67 => x"cf2ab7dc",
    68 => x"c4486e9a",
    69 => x"7258a630",
    70 => x"87c5029a",
    71 => x"c148a6c8",
    72 => x"06aac978",
    73 => x"f7c087c5",
    74 => x"c087c382",
    75 => x"66c882f0",
    76 => x"7287c702",
    77 => x"87ffc149",
    78 => x"85c184c1",
    79 => x"04adb7c8",
    80 => x"c187c7ff",
    81 => x"f0c087cf",
    82 => x"87ebc149",
    83 => x"c4c184c1",
    84 => x"7383c487",
    85 => x"6a8ac44a",
    86 => x"87f7c149",
    87 => x"4ca44970",
    88 => x"c487f2c0",
    89 => x"78c148a6",
    90 => x"c487eac0",
    91 => x"c44a7383",
    92 => x"c1496a8a",
    93 => x"84c187c1",
    94 => x"496e87db",
    95 => x"d487f8c0",
    96 => x"c0486e87",
    97 => x"c705a8e5",
    98 => x"48a6c487",
    99 => x"87c578c1",
   100 => x"e2c0496e",
   101 => x"66e0c087",
   102 => x"80c14849",
   103 => x"58a6e4c0",
   104 => x"a6c44811",
   105 => x"05987058",
   106 => x"7487cafc",
   107 => x"268ef048",
   108 => x"264c264d",
   109 => x"1e4f264b",
   110 => x"4a7186fc",
   111 => x"6949c0ff",
   112 => x"98c0c448",
   113 => x"7058a6c4",
   114 => x"87f30298",
   115 => x"fc487972",
   116 => x"0e4f268e",
   117 => x"0e5c5b5e",
   118 => x"4cc04b71",
   119 => x"029a4a13",
   120 => x"497287cd",
   121 => x"c187d0ff",
   122 => x"9a4a1384",
   123 => x"7487f305",
   124 => x"264c2648",
   125 => x"1e4f264b",
   126 => x"1e731e72",
   127 => x"02114812",
   128 => x"c34b87ca",
   129 => x"739b98df",
   130 => x"87f00288",
   131 => x"4a264b26",
   132 => x"731e4f26",
   133 => x"c11e721e",
   134 => x"87ca048b",
   135 => x"02114812",
   136 => x"028887c4",
   137 => x"4a2687f1",
   138 => x"4f264b26",
   139 => x"8148731e",
   140 => x"c502a973",
   141 => x"05531287",
   142 => x"4f2687f6",
   143 => x"711e731e",
   144 => x"4b66c84a",
   145 => x"718bc149",
   146 => x"87cf0299",
   147 => x"d4ff4812",
   148 => x"49737808",
   149 => x"99718bc1",
   150 => x"2687f105",
   151 => x"0e4f264b",
   152 => x"0e5c5b5e",
   153 => x"d4ff4a71",
   154 => x"4b66cc4c",
   155 => x"718bc149",
   156 => x"87ce0299",
   157 => x"6c7cffc3",
   158 => x"c1497352",
   159 => x"0599718b",
   160 => x"4c2687f2",
   161 => x"4f264b26",
   162 => x"ff1e731e",
   163 => x"ffc34bd4",
   164 => x"c34a6b7b",
   165 => x"496b7bff",
   166 => x"b17232c8",
   167 => x"6b7bffc3",
   168 => x"7131c84a",
   169 => x"7bffc3b2",
   170 => x"32c8496b",
   171 => x"4871b172",
   172 => x"4f264b26",
   173 => x"5c5b5e0e",
   174 => x"4d710e5d",
   175 => x"754cd4ff",
   176 => x"98ffc348",
   177 => x"e8c27c70",
   178 => x"c805bfc4",
   179 => x"4866d087",
   180 => x"a6d430c9",
   181 => x"4966d058",
   182 => x"487129d8",
   183 => x"7098ffc3",
   184 => x"4966d07c",
   185 => x"487129d0",
   186 => x"7098ffc3",
   187 => x"4966d07c",
   188 => x"487129c8",
   189 => x"7098ffc3",
   190 => x"4866d07c",
   191 => x"7098ffc3",
   192 => x"d049757c",
   193 => x"c3487129",
   194 => x"7c7098ff",
   195 => x"f0c94b6c",
   196 => x"ffc34aff",
   197 => x"87cf05ab",
   198 => x"6c7c7149",
   199 => x"028ac14b",
   200 => x"ab7187c5",
   201 => x"7387f202",
   202 => x"264d2648",
   203 => x"264b264c",
   204 => x"49c01e4f",
   205 => x"c348d4ff",
   206 => x"81c178ff",
   207 => x"a9b7c8c3",
   208 => x"2687f104",
   209 => x"5b5e0e4f",
   210 => x"c00e5d5c",
   211 => x"f7c1f0ff",
   212 => x"c0c0c14d",
   213 => x"4bc0c0c0",
   214 => x"c487d6ff",
   215 => x"c04cdff8",
   216 => x"fd49751e",
   217 => x"86c487ce",
   218 => x"c005a8c1",
   219 => x"d4ff87e5",
   220 => x"78ffc348",
   221 => x"e1c01e73",
   222 => x"49e9c1f0",
   223 => x"c487f5fc",
   224 => x"05987086",
   225 => x"d4ff87ca",
   226 => x"78ffc348",
   227 => x"87cb48c1",
   228 => x"c187defe",
   229 => x"c6ff058c",
   230 => x"2648c087",
   231 => x"264c264d",
   232 => x"0e4f264b",
   233 => x"0e5c5b5e",
   234 => x"c1f0ffc0",
   235 => x"d4ff4cc1",
   236 => x"78ffc348",
   237 => x"f849e8cf",
   238 => x"4bd387d9",
   239 => x"49741ec0",
   240 => x"c487f1fb",
   241 => x"05987086",
   242 => x"d4ff87ca",
   243 => x"78ffc348",
   244 => x"87cb48c1",
   245 => x"c187dafd",
   246 => x"dfff058b",
   247 => x"2648c087",
   248 => x"264b264c",
   249 => x"0000004f",
   250 => x"00444d43",
   251 => x"43484453",
   252 => x"69616620",
   253 => x"000a216c",
   254 => x"52524549",
   255 => x"00000000",
   256 => x"00495053",
   257 => x"74697257",
   258 => x"61662065",
   259 => x"64656c69",
   260 => x"5e0e000a",
   261 => x"0e5d5c5b",
   262 => x"ff4dffc3",
   263 => x"d0fc4bd4",
   264 => x"1eeac687",
   265 => x"c1f0e1c0",
   266 => x"c7fa49c8",
   267 => x"c186c487",
   268 => x"87c802a8",
   269 => x"c087ecfd",
   270 => x"87e8c148",
   271 => x"7087c9f9",
   272 => x"ffffcf49",
   273 => x"a9eac699",
   274 => x"fd87c802",
   275 => x"48c087d5",
   276 => x"7587d1c1",
   277 => x"4cf1c07b",
   278 => x"7087eafb",
   279 => x"ecc00298",
   280 => x"c01ec087",
   281 => x"fac1f0ff",
   282 => x"87c8f949",
   283 => x"987086c4",
   284 => x"7587da05",
   285 => x"75496b7b",
   286 => x"757b757b",
   287 => x"c17b757b",
   288 => x"c40299c0",
   289 => x"db48c187",
   290 => x"d748c087",
   291 => x"05acc287",
   292 => x"eccf87ca",
   293 => x"87fbf449",
   294 => x"87c848c0",
   295 => x"fe058cc1",
   296 => x"48c087f6",
   297 => x"4c264d26",
   298 => x"4f264b26",
   299 => x"5c5b5e0e",
   300 => x"d0ff0e5d",
   301 => x"d0e5c04d",
   302 => x"c24cc0c1",
   303 => x"c148c4e8",
   304 => x"49c0d078",
   305 => x"c787ccf4",
   306 => x"f97dc24b",
   307 => x"7dc387e3",
   308 => x"49741ec0",
   309 => x"c487ddf7",
   310 => x"05a8c186",
   311 => x"c24b87c1",
   312 => x"87cb05ab",
   313 => x"f349f8cf",
   314 => x"48c087e9",
   315 => x"c187f6c0",
   316 => x"d4ff058b",
   317 => x"87dafc87",
   318 => x"58c8e8c2",
   319 => x"cd059870",
   320 => x"c01ec187",
   321 => x"d0c1f0ff",
   322 => x"87e8f649",
   323 => x"d4ff86c4",
   324 => x"78ffc348",
   325 => x"c287eec4",
   326 => x"c258cce8",
   327 => x"48d4ff7d",
   328 => x"c178ffc3",
   329 => x"264d2648",
   330 => x"264b264c",
   331 => x"5b5e0e4f",
   332 => x"710e5d5c",
   333 => x"4cffc34d",
   334 => x"744bd4ff",
   335 => x"48d0ff7b",
   336 => x"7478c3c4",
   337 => x"c01e757b",
   338 => x"d8c1f0ff",
   339 => x"87e4f549",
   340 => x"987086c4",
   341 => x"d087cb02",
   342 => x"f6f149c4",
   343 => x"c048c187",
   344 => x"7b7487ee",
   345 => x"c87bfec3",
   346 => x"66d41ec0",
   347 => x"87ccf349",
   348 => x"7b7486c4",
   349 => x"7b747b74",
   350 => x"4ae0dad8",
   351 => x"056b7b74",
   352 => x"8ac187c5",
   353 => x"7487f505",
   354 => x"48d0ff7b",
   355 => x"48c078c2",
   356 => x"4c264d26",
   357 => x"4f264b26",
   358 => x"5c5b5e0e",
   359 => x"86fc0e5d",
   360 => x"d4ff4b71",
   361 => x"c57ec04c",
   362 => x"4adfcdee",
   363 => x"6c7cffc3",
   364 => x"a8fec348",
   365 => x"87f8c005",
   366 => x"9b734d74",
   367 => x"d487cc02",
   368 => x"49731e66",
   369 => x"c487d8f2",
   370 => x"ff87d486",
   371 => x"d1c448d0",
   372 => x"4a66d478",
   373 => x"c17dffc3",
   374 => x"87f8058a",
   375 => x"c35aa6d8",
   376 => x"737c7cff",
   377 => x"87c5059b",
   378 => x"d048d0ff",
   379 => x"7e4ac178",
   380 => x"fe058ac1",
   381 => x"486e87f6",
   382 => x"4d268efc",
   383 => x"4b264c26",
   384 => x"731e4f26",
   385 => x"c04a711e",
   386 => x"48d4ff4b",
   387 => x"ff78ffc3",
   388 => x"c3c448d0",
   389 => x"48d4ff78",
   390 => x"7278ffc3",
   391 => x"f0ffc01e",
   392 => x"f249d1c1",
   393 => x"86c487ce",
   394 => x"d2059870",
   395 => x"1ec0c887",
   396 => x"fd4966cc",
   397 => x"86c487e2",
   398 => x"d0ff4b70",
   399 => x"7378c248",
   400 => x"264b2648",
   401 => x"5b5e0e4f",
   402 => x"c00e5d5c",
   403 => x"f0ffc01e",
   404 => x"f149c9c1",
   405 => x"1ed287de",
   406 => x"49d4e8c2",
   407 => x"c887f9fc",
   408 => x"c14cc086",
   409 => x"acb7d284",
   410 => x"c287f804",
   411 => x"bf97d4e8",
   412 => x"99c0c349",
   413 => x"05a9c0c1",
   414 => x"c287e7c0",
   415 => x"bf97dbe8",
   416 => x"c231d049",
   417 => x"bf97dce8",
   418 => x"7232c84a",
   419 => x"dde8c2b1",
   420 => x"b14abf97",
   421 => x"ffcf4c71",
   422 => x"c19cffff",
   423 => x"c134ca84",
   424 => x"e8c287e7",
   425 => x"49bf97dd",
   426 => x"99c631c1",
   427 => x"97dee8c2",
   428 => x"b7c74abf",
   429 => x"c2b1722a",
   430 => x"bf97d9e8",
   431 => x"9dcf4d4a",
   432 => x"97dae8c2",
   433 => x"9ac34abf",
   434 => x"e8c232ca",
   435 => x"4bbf97db",
   436 => x"b27333c2",
   437 => x"97dce8c2",
   438 => x"c0c34bbf",
   439 => x"2bb7c69b",
   440 => x"81c2b273",
   441 => x"307148c1",
   442 => x"48c14970",
   443 => x"4d703075",
   444 => x"84c14c72",
   445 => x"c0c89471",
   446 => x"cc06adb7",
   447 => x"b734c187",
   448 => x"b7c0c82d",
   449 => x"f4ff01ad",
   450 => x"26487487",
   451 => x"264c264d",
   452 => x"0e4f264b",
   453 => x"5d5c5b5e",
   454 => x"c286fc0e",
   455 => x"c048fcf0",
   456 => x"f4e8c278",
   457 => x"fb49c01e",
   458 => x"86c487d8",
   459 => x"c5059870",
   460 => x"c948c087",
   461 => x"4dc087d7",
   462 => x"48f8f5c2",
   463 => x"e9c278c1",
   464 => x"e6c04aea",
   465 => x"4bc849e4",
   466 => x"7087c7eb",
   467 => x"87c60598",
   468 => x"48f8f5c2",
   469 => x"eac278c0",
   470 => x"e6c04ac6",
   471 => x"4bc849f0",
   472 => x"7087efea",
   473 => x"87c60598",
   474 => x"48f8f5c2",
   475 => x"f5c278c0",
   476 => x"c002bff8",
   477 => x"efc287ff",
   478 => x"c24dbffa",
   479 => x"bf9ff2f0",
   480 => x"58a6c448",
   481 => x"a8ead6c5",
   482 => x"c287c705",
   483 => x"4dbffaef",
   484 => x"486e87ce",
   485 => x"a8d5e9ca",
   486 => x"c087c502",
   487 => x"87edc748",
   488 => x"1ef4e8c2",
   489 => x"d9f94975",
   490 => x"7086c487",
   491 => x"87c50598",
   492 => x"d8c748c0",
   493 => x"c6eac287",
   494 => x"fce6c04a",
   495 => x"e94bc849",
   496 => x"987087d0",
   497 => x"87c8c005",
   498 => x"48fcf0c2",
   499 => x"87d878c1",
   500 => x"4aeae9c2",
   501 => x"49c8e7c0",
   502 => x"f5e84bc8",
   503 => x"02987087",
   504 => x"c087c5c0",
   505 => x"87e5c648",
   506 => x"97f2f0c2",
   507 => x"d5c149bf",
   508 => x"cdc005a9",
   509 => x"f3f0c287",
   510 => x"c249bf97",
   511 => x"c002a9ea",
   512 => x"48c087c5",
   513 => x"c287c6c6",
   514 => x"bf97f4e8",
   515 => x"58a6c448",
   516 => x"02a8e9c3",
   517 => x"6e87cec0",
   518 => x"a8ebc348",
   519 => x"87c5c002",
   520 => x"e8c548c0",
   521 => x"ffe8c287",
   522 => x"9949bf97",
   523 => x"87ccc005",
   524 => x"97c0e9c2",
   525 => x"a9c249bf",
   526 => x"87c5c002",
   527 => x"ccc548c0",
   528 => x"c1e9c287",
   529 => x"c248bf97",
   530 => x"7058f8f0",
   531 => x"88c1484c",
   532 => x"58fcf0c2",
   533 => x"97c2e9c2",
   534 => x"817549bf",
   535 => x"97c3e9c2",
   536 => x"32c84abf",
   537 => x"c27ea172",
   538 => x"6e48d4f5",
   539 => x"c4e9c278",
   540 => x"c248bf97",
   541 => x"c258ecf5",
   542 => x"02bffcf0",
   543 => x"c287d3c2",
   544 => x"c04ac6ea",
   545 => x"c849d8e6",
   546 => x"87c6e64b",
   547 => x"c0029870",
   548 => x"48c087c5",
   549 => x"c287f6c3",
   550 => x"4cbff4f0",
   551 => x"5ce8f5c2",
   552 => x"97d9e9c2",
   553 => x"31c849bf",
   554 => x"97d8e9c2",
   555 => x"49a14abf",
   556 => x"97dae9c2",
   557 => x"32d04abf",
   558 => x"c249a172",
   559 => x"bf97dbe9",
   560 => x"7232d84a",
   561 => x"f5c249a1",
   562 => x"f5c259f0",
   563 => x"c291bfe8",
   564 => x"81bfd4f5",
   565 => x"59dcf5c2",
   566 => x"97e1e9c2",
   567 => x"32c84abf",
   568 => x"97e0e9c2",
   569 => x"4aa24bbf",
   570 => x"97e2e9c2",
   571 => x"33d04bbf",
   572 => x"c24aa273",
   573 => x"bf97e3e9",
   574 => x"d89bcf4b",
   575 => x"4aa27333",
   576 => x"5ae0f5c2",
   577 => x"92748ac2",
   578 => x"48e0f5c2",
   579 => x"c178a172",
   580 => x"e9c287c7",
   581 => x"49bf97c6",
   582 => x"e9c231c8",
   583 => x"4abf97c5",
   584 => x"31c549a1",
   585 => x"c981ffc7",
   586 => x"e8f5c229",
   587 => x"cbe9c259",
   588 => x"c84abf97",
   589 => x"cae9c232",
   590 => x"a24bbf97",
   591 => x"f0f5c24a",
   592 => x"e8f5c25a",
   593 => x"826e92bf",
   594 => x"5ae4f5c2",
   595 => x"48dcf5c2",
   596 => x"f5c278c0",
   597 => x"a17248d8",
   598 => x"f0f5c278",
   599 => x"dcf5c248",
   600 => x"f5c278bf",
   601 => x"f5c248f4",
   602 => x"c278bfe0",
   603 => x"02bffcf0",
   604 => x"7487c9c0",
   605 => x"a630c448",
   606 => x"87c9c058",
   607 => x"bfe4f5c2",
   608 => x"a630c448",
   609 => x"c0f1c258",
   610 => x"c1786e48",
   611 => x"268efc48",
   612 => x"264c264d",
   613 => x"004f264b",
   614 => x"33544146",
   615 => x"20202032",
   616 => x"00000000",
   617 => x"31544146",
   618 => x"20202036",
   619 => x"00000000",
   620 => x"33544146",
   621 => x"20202032",
   622 => x"00000000",
   623 => x"33544146",
   624 => x"20202032",
   625 => x"00000000",
   626 => x"31544146",
   627 => x"20202036",
   628 => x"5b5e0e00",
   629 => x"710e5d5c",
   630 => x"fcf0c24a",
   631 => x"87cb02bf",
   632 => x"2bc74b72",
   633 => x"ffc14d72",
   634 => x"7287c99d",
   635 => x"722bc84b",
   636 => x"9dffc34d",
   637 => x"bfd4f5c2",
   638 => x"dcfec083",
   639 => x"d902abbf",
   640 => x"e0fec087",
   641 => x"f4e8c25b",
   642 => x"ef49731e",
   643 => x"86c487f4",
   644 => x"c5059870",
   645 => x"c048c087",
   646 => x"f0c287e6",
   647 => x"d202bffc",
   648 => x"c4497587",
   649 => x"f4e8c291",
   650 => x"cf4c6981",
   651 => x"ffffffff",
   652 => x"7587cb9c",
   653 => x"c291c249",
   654 => x"9f81f4e8",
   655 => x"48744c69",
   656 => x"4c264d26",
   657 => x"4f264b26",
   658 => x"5c5b5e0e",
   659 => x"86f40e5d",
   660 => x"c459a6c8",
   661 => x"80c84866",
   662 => x"6e58a6c4",
   663 => x"1e78c048",
   664 => x"ffcc49c1",
   665 => x"7086c487",
   666 => x"c0029c4c",
   667 => x"f1c287fc",
   668 => x"66dc4ac4",
   669 => x"feddff49",
   670 => x"02987087",
   671 => x"7487ebc0",
   672 => x"4966dc4a",
   673 => x"deff4bcb",
   674 => x"987087c8",
   675 => x"c087db02",
   676 => x"029c741e",
   677 => x"4dc087c4",
   678 => x"4dc187c2",
   679 => x"c3cc4975",
   680 => x"7086c487",
   681 => x"ff059c4c",
   682 => x"9c7487c4",
   683 => x"87f5c102",
   684 => x"6e49a4dc",
   685 => x"da786948",
   686 => x"66c449a4",
   687 => x"9f85c44d",
   688 => x"f0c27d69",
   689 => x"d302bffc",
   690 => x"49a4d487",
   691 => x"c049699f",
   692 => x"7199ffff",
   693 => x"c430d048",
   694 => x"87c258a6",
   695 => x"496e7ec0",
   696 => x"70806d48",
   697 => x"4866c47d",
   698 => x"66c478c0",
   699 => x"6d81cc49",
   700 => x"4966c479",
   701 => x"79c081d0",
   702 => x"c048a6c8",
   703 => x"4c66c878",
   704 => x"d44a66c4",
   705 => x"c8497482",
   706 => x"49a17291",
   707 => x"796d41c0",
   708 => x"b7c684c1",
   709 => x"e7ff04ac",
   710 => x"4966c487",
   711 => x"c081c4c1",
   712 => x"c248c179",
   713 => x"f448c087",
   714 => x"264d268e",
   715 => x"264b264c",
   716 => x"5b5e0e4f",
   717 => x"710e5d5c",
   718 => x"4d66d04c",
   719 => x"7585496c",
   720 => x"f8f0c2b9",
   721 => x"baff4abf",
   722 => x"99719972",
   723 => x"87e4c002",
   724 => x"6b4ba4c4",
   725 => x"87f9f949",
   726 => x"f0c27b70",
   727 => x"6c49bff4",
   728 => x"757c7181",
   729 => x"f8f0c2b9",
   730 => x"baff4abf",
   731 => x"99719972",
   732 => x"87dcff05",
   733 => x"4d267c75",
   734 => x"4b264c26",
   735 => x"731e4f26",
   736 => x"c24b711e",
   737 => x"49bfd8f5",
   738 => x"6a4aa3c4",
   739 => x"c28ac24a",
   740 => x"92bff4f0",
   741 => x"c249a172",
   742 => x"4abff8f0",
   743 => x"a1729a6b",
   744 => x"e0fec049",
   745 => x"1e66c859",
   746 => x"87d6e971",
   747 => x"987086c4",
   748 => x"c087c405",
   749 => x"c187c248",
   750 => x"264b2648",
   751 => x"1e731e4f",
   752 => x"f5c24b71",
   753 => x"c449bfd8",
   754 => x"4a6a4aa3",
   755 => x"f0c28ac2",
   756 => x"7292bff4",
   757 => x"f0c249a1",
   758 => x"6b4abff8",
   759 => x"49a1729a",
   760 => x"59e0fec0",
   761 => x"711e66c8",
   762 => x"c487c2e5",
   763 => x"05987086",
   764 => x"48c087c4",
   765 => x"48c187c2",
   766 => x"4f264b26",
   767 => x"5c5b5e0e",
   768 => x"86e40e5d",
   769 => x"ecc04b71",
   770 => x"28c94866",
   771 => x"c258a6cc",
   772 => x"49bff8f0",
   773 => x"4871b9ff",
   774 => x"d49866c8",
   775 => x"487158a6",
   776 => x"a6d0986b",
   777 => x"7ea3c458",
   778 => x"6e48a6c4",
   779 => x"66d078bf",
   780 => x"a866cc48",
   781 => x"c887c605",
   782 => x"c7c37b66",
   783 => x"48a6d487",
   784 => x"ffffffc1",
   785 => x"c478ffff",
   786 => x"c078ff80",
   787 => x"4da3d44a",
   788 => x"91c84972",
   789 => x"d049a175",
   790 => x"8c694c66",
   791 => x"04acb7c0",
   792 => x"66d487cd",
   793 => x"c603acb7",
   794 => x"5aa6dc87",
   795 => x"c15ca6d8",
   796 => x"aab7c682",
   797 => x"87d5ff04",
   798 => x"c04866d8",
   799 => x"d004a8b7",
   800 => x"4966d887",
   801 => x"a17591c8",
   802 => x"6e7b2149",
   803 => x"c9786948",
   804 => x"cc7bc087",
   805 => x"486e49a3",
   806 => x"66c87869",
   807 => x"cc886b48",
   808 => x"f0c258a6",
   809 => x"c848bff4",
   810 => x"58a6c490",
   811 => x"6e4866c8",
   812 => x"87c901a8",
   813 => x"6e4866c8",
   814 => x"fdc003a8",
   815 => x"a3c4c187",
   816 => x"49bf6e7e",
   817 => x"a17591c8",
   818 => x"7966cc49",
   819 => x"c849bf6e",
   820 => x"49a17591",
   821 => x"796681c4",
   822 => x"6e48a6d0",
   823 => x"66d078bf",
   824 => x"05a8c548",
   825 => x"a6c487c7",
   826 => x"c878c048",
   827 => x"4866d087",
   828 => x"a6c880c1",
   829 => x"c4486e58",
   830 => x"66c87866",
   831 => x"f849731e",
   832 => x"86c487ef",
   833 => x"1ef4e8c2",
   834 => x"f1f94973",
   835 => x"49a3d087",
   836 => x"7966f0c0",
   837 => x"4d268ee0",
   838 => x"4b264c26",
   839 => x"5e0e4f26",
   840 => x"710e5c5b",
   841 => x"724bc04a",
   842 => x"e0c0029a",
   843 => x"49a2da87",
   844 => x"c24b699f",
   845 => x"02bffcf0",
   846 => x"a2d487cf",
   847 => x"49699f49",
   848 => x"ffffc04c",
   849 => x"c234d09c",
   850 => x"744cc087",
   851 => x"029b73b3",
   852 => x"c24a87df",
   853 => x"f4f0c28a",
   854 => x"c29249bf",
   855 => x"48bfd8f5",
   856 => x"f5c28072",
   857 => x"487158f8",
   858 => x"f1c230c4",
   859 => x"e9c058c4",
   860 => x"dcf5c287",
   861 => x"f5c24bbf",
   862 => x"f5c248f4",
   863 => x"c278bfe0",
   864 => x"02bffcf0",
   865 => x"f0c287c9",
   866 => x"c449bff4",
   867 => x"c287c731",
   868 => x"49bfe4f5",
   869 => x"f1c231c4",
   870 => x"f5c259c4",
   871 => x"4c265bf4",
   872 => x"4f264b26",
   873 => x"5c5b5e0e",
   874 => x"86f00e5d",
   875 => x"cf59a6c8",
   876 => x"f8ffffff",
   877 => x"c47ec04c",
   878 => x"87d80266",
   879 => x"48f0e8c2",
   880 => x"e8c278c0",
   881 => x"f5c248e8",
   882 => x"c278bff4",
   883 => x"c248ece8",
   884 => x"78bff0f5",
   885 => x"48d1f1c2",
   886 => x"f1c250c0",
   887 => x"c249bfc0",
   888 => x"4abff0e8",
   889 => x"c403aa71",
   890 => x"497287cc",
   891 => x"c00599cf",
   892 => x"fec087ea",
   893 => x"e8c248dc",
   894 => x"c278bfe8",
   895 => x"c21ef4e8",
   896 => x"49bfe8e8",
   897 => x"48e8e8c2",
   898 => x"7178a1c1",
   899 => x"87f2dfff",
   900 => x"fec086c4",
   901 => x"e8c248d8",
   902 => x"87cc78f4",
   903 => x"bfd8fec0",
   904 => x"80e0c048",
   905 => x"58dcfec0",
   906 => x"bff0e8c2",
   907 => x"c280c148",
   908 => x"2758f4e8",
   909 => x"00000f98",
   910 => x"4dbf97bf",
   911 => x"e5c2029d",
   912 => x"ade5c387",
   913 => x"87dec202",
   914 => x"bfd8fec0",
   915 => x"49a3cb4b",
   916 => x"accf4c11",
   917 => x"87d2c105",
   918 => x"99df4975",
   919 => x"91cd89c1",
   920 => x"81c4f1c2",
   921 => x"124aa3c1",
   922 => x"4aa3c351",
   923 => x"a3c55112",
   924 => x"c751124a",
   925 => x"51124aa3",
   926 => x"124aa3c9",
   927 => x"4aa3ce51",
   928 => x"a3d05112",
   929 => x"d251124a",
   930 => x"51124aa3",
   931 => x"124aa3d4",
   932 => x"4aa3d651",
   933 => x"a3d85112",
   934 => x"dc51124a",
   935 => x"51124aa3",
   936 => x"124aa3de",
   937 => x"c07ec151",
   938 => x"497487fc",
   939 => x"c00599c8",
   940 => x"497487ed",
   941 => x"d30599d0",
   942 => x"66e0c087",
   943 => x"87ccc002",
   944 => x"e0c04973",
   945 => x"98700f66",
   946 => x"87d3c002",
   947 => x"c6c0056e",
   948 => x"c4f1c287",
   949 => x"c050c048",
   950 => x"48bfd8fe",
   951 => x"c287e9c2",
   952 => x"c048d1f1",
   953 => x"f1c27e50",
   954 => x"c249bfc0",
   955 => x"4abff0e8",
   956 => x"fb04aa71",
   957 => x"ffcf87f4",
   958 => x"4cf8ffff",
   959 => x"bff4f5c2",
   960 => x"87c8c005",
   961 => x"bffcf0c2",
   962 => x"87fac102",
   963 => x"bfece8c2",
   964 => x"87fdea49",
   965 => x"58f0e8c2",
   966 => x"c248a6c4",
   967 => x"78bfece8",
   968 => x"bffcf0c2",
   969 => x"87dbc002",
   970 => x"744966c4",
   971 => x"02a97499",
   972 => x"c887c8c0",
   973 => x"78c048a6",
   974 => x"c887e7c0",
   975 => x"78c148a6",
   976 => x"c487dfc0",
   977 => x"ffcf4966",
   978 => x"02a999f8",
   979 => x"cc87c8c0",
   980 => x"78c048a6",
   981 => x"cc87c5c0",
   982 => x"78c148a6",
   983 => x"cc48a6c8",
   984 => x"66c87866",
   985 => x"87dec005",
   986 => x"c24966c4",
   987 => x"f4f0c289",
   988 => x"f5c291bf",
   989 => x"7148bfd8",
   990 => x"ece8c280",
   991 => x"f0e8c258",
   992 => x"f978c048",
   993 => x"48c087d4",
   994 => x"ffffffcf",
   995 => x"8ef04cf8",
   996 => x"4c264d26",
   997 => x"4f264b26",
   998 => x"00000000",
   999 => x"ffffffff",
  1000 => x"48d4ff1e",
  1001 => x"6878ffc3",
  1002 => x"1e4f2648",
  1003 => x"c348d4ff",
  1004 => x"d0ff78ff",
  1005 => x"78e1c048",
  1006 => x"d448d4ff",
  1007 => x"1e4f2678",
  1008 => x"c048d0ff",
  1009 => x"4f2678e0",
  1010 => x"87d4ff1e",
  1011 => x"02994970",
  1012 => x"fbc087c6",
  1013 => x"87f105a9",
  1014 => x"4f264871",
  1015 => x"5c5b5e0e",
  1016 => x"c04b710e",
  1017 => x"87f8fe4c",
  1018 => x"02994970",
  1019 => x"c087f9c0",
  1020 => x"c002a9ec",
  1021 => x"fbc087f2",
  1022 => x"ebc002a9",
  1023 => x"b766cc87",
  1024 => x"87c703ac",
  1025 => x"c20266d0",
  1026 => x"71537187",
  1027 => x"87c20299",
  1028 => x"cbfe84c1",
  1029 => x"99497087",
  1030 => x"c087cd02",
  1031 => x"c702a9ec",
  1032 => x"a9fbc087",
  1033 => x"87d5ff05",
  1034 => x"c30266d0",
  1035 => x"7b97c087",
  1036 => x"05a9fbc0",
  1037 => x"4a7487c7",
  1038 => x"c28a0ac0",
  1039 => x"724a7487",
  1040 => x"264c2648",
  1041 => x"1e4f264b",
  1042 => x"7087d5fd",
  1043 => x"a9f0c049",
  1044 => x"c087c904",
  1045 => x"c301a9f9",
  1046 => x"89f0c087",
  1047 => x"04a9c1c1",
  1048 => x"dac187c9",
  1049 => x"87c301a9",
  1050 => x"7189f7c0",
  1051 => x"0e4f2648",
  1052 => x"5d5c5b5e",
  1053 => x"7186f80e",
  1054 => x"fc7ec04c",
  1055 => x"4bc087ed",
  1056 => x"97d0c4c1",
  1057 => x"a9c049bf",
  1058 => x"fc87cf04",
  1059 => x"83c187fa",
  1060 => x"97d0c4c1",
  1061 => x"06ab49bf",
  1062 => x"c4c187f1",
  1063 => x"02bf97d0",
  1064 => x"fbfb87cf",
  1065 => x"99497087",
  1066 => x"c087c602",
  1067 => x"f105a9ec",
  1068 => x"fb4bc087",
  1069 => x"4d7087ea",
  1070 => x"c887e5fb",
  1071 => x"dffb58a6",
  1072 => x"c14a7087",
  1073 => x"49a4c883",
  1074 => x"ad496997",
  1075 => x"c987da05",
  1076 => x"699749a4",
  1077 => x"a966c449",
  1078 => x"ca87ce05",
  1079 => x"699749a4",
  1080 => x"c405aa49",
  1081 => x"d07ec187",
  1082 => x"adecc087",
  1083 => x"c087c602",
  1084 => x"c405adfb",
  1085 => x"c14bc087",
  1086 => x"fe026e7e",
  1087 => x"fefa87f5",
  1088 => x"f8487387",
  1089 => x"264d268e",
  1090 => x"264b264c",
  1091 => x"0000004f",
  1092 => x"1e731e00",
  1093 => x"c84bd4ff",
  1094 => x"d0ff4a66",
  1095 => x"78c5c848",
  1096 => x"c148d4ff",
  1097 => x"7b1178d4",
  1098 => x"f9058ac1",
  1099 => x"48d0ff87",
  1100 => x"4b2678c4",
  1101 => x"5e0e4f26",
  1102 => x"0e5d5c5b",
  1103 => x"a6c486f8",
  1104 => x"c21e6e59",
  1105 => x"e349c8f6",
  1106 => x"86c487fe",
  1107 => x"c4029870",
  1108 => x"f2c187ee",
  1109 => x"6e4cbfc8",
  1110 => x"87d3fc49",
  1111 => x"c158a6c8",
  1112 => x"fe1eccca",
  1113 => x"c487e5fc",
  1114 => x"c5056686",
  1115 => x"48a6c487",
  1116 => x"d0ff78c1",
  1117 => x"ff78c548",
  1118 => x"d5c148d4",
  1119 => x"4966c478",
  1120 => x"31c689c1",
  1121 => x"97c0f2c1",
  1122 => x"71484abf",
  1123 => x"08d4ffb0",
  1124 => x"48d0ff78",
  1125 => x"f6c278c4",
  1126 => x"49bf97c4",
  1127 => x"dd0299d0",
  1128 => x"ff78c587",
  1129 => x"d6c148d4",
  1130 => x"ff4ac078",
  1131 => x"ffc348d4",
  1132 => x"c082c178",
  1133 => x"f204aae0",
  1134 => x"48d0ff87",
  1135 => x"d4ff78c4",
  1136 => x"78ffc348",
  1137 => x"c548d0ff",
  1138 => x"48d4ff78",
  1139 => x"c178d3c1",
  1140 => x"48d0ff78",
  1141 => x"b7c078c4",
  1142 => x"ccc206ac",
  1143 => x"d0f6c287",
  1144 => x"c48c4bbf",
  1145 => x"9b735ca6",
  1146 => x"87ddc102",
  1147 => x"8b4dc0c8",
  1148 => x"03abb7c0",
  1149 => x"c0c887c6",
  1150 => x"4bc04da3",
  1151 => x"97c4f6c2",
  1152 => x"99d049bf",
  1153 => x"c087cf02",
  1154 => x"c8f6c21e",
  1155 => x"87eee549",
  1156 => x"4c7086c4",
  1157 => x"e8c287d8",
  1158 => x"f6c21ef4",
  1159 => x"dde549c8",
  1160 => x"754c7087",
  1161 => x"f4e8c21e",
  1162 => x"87e5fb49",
  1163 => x"9c7486c8",
  1164 => x"c087c505",
  1165 => x"87cac148",
  1166 => x"f6c21ec1",
  1167 => x"f0e349c8",
  1168 => x"7386c487",
  1169 => x"e3fe059b",
  1170 => x"c04c6e87",
  1171 => x"d106acb7",
  1172 => x"c8f6c287",
  1173 => x"d078c048",
  1174 => x"f478c080",
  1175 => x"d4f6c280",
  1176 => x"b7c078bf",
  1177 => x"f4fd01ac",
  1178 => x"48d0ff87",
  1179 => x"d4ff78c5",
  1180 => x"78d3c148",
  1181 => x"d0ff78c0",
  1182 => x"c178c448",
  1183 => x"87c2c048",
  1184 => x"8ef848c0",
  1185 => x"4c264d26",
  1186 => x"4f264b26",
  1187 => x"20746f47",
  1188 => x"69747865",
  1189 => x"0000646e",
  1190 => x"64616f4c",
  1191 => x"2e676e69",
  1192 => x"00002e2e",
  1193 => x"61422080",
  1194 => x"00006b63",
  1195 => x"64616f4c",
  1196 => x"202e2a20",
  1197 => x"00000000",
  1198 => x"0000203a",
  1199 => x"61422080",
  1200 => x"00006b63",
  1201 => x"78452080",
  1202 => x"00007469",
  1203 => x"49204453",
  1204 => x"2e74696e",
  1205 => x"0000002e",
  1206 => x"00004b4f",
  1207 => x"544f4f42",
  1208 => x"20202020",
  1209 => x"004d4f52",
  1210 => x"5c5b5e0e",
  1211 => x"86fc0e5d",
  1212 => x"4bc04d71",
  1213 => x"c004ad4c",
  1214 => x"c1c187e8",
  1215 => x"9c741eef",
  1216 => x"c087c402",
  1217 => x"c187c24a",
  1218 => x"ea49724a",
  1219 => x"86c487d6",
  1220 => x"83c158a6",
  1221 => x"87c2056e",
  1222 => x"84c14b75",
  1223 => x"ff06ab75",
  1224 => x"486e87d8",
  1225 => x"4d268efc",
  1226 => x"4b264c26",
  1227 => x"5e0e4f26",
  1228 => x"710e5c5b",
  1229 => x"0266cc4b",
  1230 => x"c04c87d8",
  1231 => x"d8028cf0",
  1232 => x"c14a7487",
  1233 => x"87d1028a",
  1234 => x"87cd028a",
  1235 => x"87c9028a",
  1236 => x"497387d9",
  1237 => x"d287dff7",
  1238 => x"c01e7487",
  1239 => x"f9d7c149",
  1240 => x"731e7487",
  1241 => x"f1d7c149",
  1242 => x"2686c887",
  1243 => x"264b264c",
  1244 => x"5b5e0e4f",
  1245 => x"fc0e5d5c",
  1246 => x"494c7186",
  1247 => x"f7c291de",
  1248 => x"85714de8",
  1249 => x"c1026d97",
  1250 => x"f7c287db",
  1251 => x"7449bfd8",
  1252 => x"d3fd7181",
  1253 => x"58a6c487",
  1254 => x"f2c0026e",
  1255 => x"dcf7c287",
  1256 => x"cb4a6e4b",
  1257 => x"c3fafe49",
  1258 => x"cc4b7487",
  1259 => x"ccf2c193",
  1260 => x"c183c483",
  1261 => x"747bd8ca",
  1262 => x"dfc1c149",
  1263 => x"c17b7587",
  1264 => x"bf97c4f2",
  1265 => x"f7c21e49",
  1266 => x"e1fd49dc",
  1267 => x"7486c487",
  1268 => x"c7c1c149",
  1269 => x"c149c087",
  1270 => x"c287e3c2",
  1271 => x"c048c0f6",
  1272 => x"eddf4950",
  1273 => x"268efc87",
  1274 => x"264c264d",
  1275 => x"1e4f264b",
  1276 => x"4b711e73",
  1277 => x"d8f7c249",
  1278 => x"fb7181bf",
  1279 => x"4a7087ea",
  1280 => x"87c4029a",
  1281 => x"87d6e449",
  1282 => x"48d8f7c2",
  1283 => x"497378c0",
  1284 => x"2687fac1",
  1285 => x"1e4f264b",
  1286 => x"4b711e73",
  1287 => x"024aa3c4",
  1288 => x"c187d0c1",
  1289 => x"87dc028a",
  1290 => x"f2c0028a",
  1291 => x"c1058a87",
  1292 => x"f7c287d3",
  1293 => x"c102bfd8",
  1294 => x"c14887cb",
  1295 => x"dcf7c288",
  1296 => x"87c1c158",
  1297 => x"bfd8f7c2",
  1298 => x"c289c649",
  1299 => x"c059dcf7",
  1300 => x"c003a9b7",
  1301 => x"f7c287ef",
  1302 => x"78c048d8",
  1303 => x"c287e6c0",
  1304 => x"02bfd4f7",
  1305 => x"f7c287df",
  1306 => x"c148bfd8",
  1307 => x"dcf7c280",
  1308 => x"c287d258",
  1309 => x"02bfd4f7",
  1310 => x"f7c287cb",
  1311 => x"c648bfd8",
  1312 => x"dcf7c280",
  1313 => x"c4497358",
  1314 => x"264b2687",
  1315 => x"5b5e0e4f",
  1316 => x"f00e5d5c",
  1317 => x"59a6d086",
  1318 => x"4df4e8c2",
  1319 => x"f7c24cc0",
  1320 => x"78c148d4",
  1321 => x"c048a6c8",
  1322 => x"5da6c478",
  1323 => x"bfd8f7c2",
  1324 => x"06a8c048",
  1325 => x"c887c1c1",
  1326 => x"a6c45ca6",
  1327 => x"f4e8c25d",
  1328 => x"c0029848",
  1329 => x"66c487f2",
  1330 => x"efc1c14d",
  1331 => x"0266cc1e",
  1332 => x"4cc087c4",
  1333 => x"4cc187c2",
  1334 => x"c7e34974",
  1335 => x"a686c487",
  1336 => x"c885c158",
  1337 => x"80c14866",
  1338 => x"c258a6cc",
  1339 => x"adbfd8f7",
  1340 => x"6e87c503",
  1341 => x"87d1ff05",
  1342 => x"4cc04d6e",
  1343 => x"c3029d75",
  1344 => x"c1c187db",
  1345 => x"66cc1eef",
  1346 => x"c887c702",
  1347 => x"78c048a6",
  1348 => x"a6c887c5",
  1349 => x"c878c148",
  1350 => x"c7e24966",
  1351 => x"a686c487",
  1352 => x"c2026e58",
  1353 => x"cb4987e4",
  1354 => x"49699781",
  1355 => x"c10299d0",
  1356 => x"497487d4",
  1357 => x"f2c191cc",
  1358 => x"cfc181cc",
  1359 => x"81c879ef",
  1360 => x"7451ffc3",
  1361 => x"c291de49",
  1362 => x"714de8f7",
  1363 => x"97c1c285",
  1364 => x"49a5c17d",
  1365 => x"c251e0c0",
  1366 => x"bf97c4f1",
  1367 => x"c187d202",
  1368 => x"4ba5c284",
  1369 => x"4ac4f1c2",
  1370 => x"f2fe49db",
  1371 => x"d9c187fe",
  1372 => x"49a5cd87",
  1373 => x"84c151c0",
  1374 => x"6e4ba5c2",
  1375 => x"fe49cb4a",
  1376 => x"c187e9f2",
  1377 => x"497487c4",
  1378 => x"f2c191cc",
  1379 => x"cdc181cc",
  1380 => x"f1c279f1",
  1381 => x"02bf97c4",
  1382 => x"497487d8",
  1383 => x"84c191de",
  1384 => x"4be8f7c2",
  1385 => x"f1c28371",
  1386 => x"49dd4ac4",
  1387 => x"87fcf1fe",
  1388 => x"4b7487d8",
  1389 => x"f7c293de",
  1390 => x"a3cb83e8",
  1391 => x"c151c049",
  1392 => x"4a6e7384",
  1393 => x"f1fe49cb",
  1394 => x"66c887e2",
  1395 => x"cc80c148",
  1396 => x"acc758a6",
  1397 => x"87c5c003",
  1398 => x"e5fc056e",
  1399 => x"03acc787",
  1400 => x"c287e4c0",
  1401 => x"c048d4f7",
  1402 => x"cc497478",
  1403 => x"ccf2c191",
  1404 => x"f1cdc181",
  1405 => x"de497479",
  1406 => x"e8f7c291",
  1407 => x"c151c081",
  1408 => x"04acc784",
  1409 => x"c187dcff",
  1410 => x"c048e8f3",
  1411 => x"e0f3c150",
  1412 => x"ead9c148",
  1413 => x"c180c478",
  1414 => x"c878e4ca",
  1415 => x"d7d0c180",
  1416 => x"4966cc78",
  1417 => x"87f4f7c0",
  1418 => x"4d268ef0",
  1419 => x"4b264c26",
  1420 => x"731e4f26",
  1421 => x"494b711e",
  1422 => x"f2c191cc",
  1423 => x"a1c881cc",
  1424 => x"c0f2c14a",
  1425 => x"c9501248",
  1426 => x"c4c14aa1",
  1427 => x"501248d0",
  1428 => x"f2c181ca",
  1429 => x"501148c4",
  1430 => x"f0f84973",
  1431 => x"264b2687",
  1432 => x"49c01e4f",
  1433 => x"87d6f8c0",
  1434 => x"711e4f26",
  1435 => x"91cc494a",
  1436 => x"81ccf2c1",
  1437 => x"f6c281c8",
  1438 => x"501148c0",
  1439 => x"49a2f0c0",
  1440 => x"87f3ecfe",
  1441 => x"c9d549c0",
  1442 => x"1e4f2687",
  1443 => x"c34ad4ff",
  1444 => x"d0ff7aff",
  1445 => x"78e1c048",
  1446 => x"7a717ade",
  1447 => x"28b7c848",
  1448 => x"48717a70",
  1449 => x"7028b7d0",
  1450 => x"d848717a",
  1451 => x"7a7028b7",
  1452 => x"c048d0ff",
  1453 => x"4f2678e0",
  1454 => x"5c5b5e0e",
  1455 => x"86f40e5d",
  1456 => x"cc494d71",
  1457 => x"ccf2c191",
  1458 => x"4aa1c881",
  1459 => x"c47ea1ca",
  1460 => x"f5c248a6",
  1461 => x"6e78bffc",
  1462 => x"c44bbf97",
  1463 => x"2c734c66",
  1464 => x"a6cc4812",
  1465 => x"c19c7058",
  1466 => x"9781c984",
  1467 => x"acb74969",
  1468 => x"c087c204",
  1469 => x"bf976e4c",
  1470 => x"4966c84a",
  1471 => x"b9ff3172",
  1472 => x"749966c4",
  1473 => x"70307248",
  1474 => x"f6c2b14a",
  1475 => x"fd7159c0",
  1476 => x"1ec787f9",
  1477 => x"bfd0f7c2",
  1478 => x"ccf2c11e",
  1479 => x"c0f6c21e",
  1480 => x"c149bf97",
  1481 => x"497587f4",
  1482 => x"87f0f3c0",
  1483 => x"4d268ee8",
  1484 => x"4b264c26",
  1485 => x"731e4f26",
  1486 => x"494b711e",
  1487 => x"7387f9fd",
  1488 => x"87f4fd49",
  1489 => x"4f264b26",
  1490 => x"711e731e",
  1491 => x"4aa3c24b",
  1492 => x"c187d602",
  1493 => x"e2c0058a",
  1494 => x"d0f7c287",
  1495 => x"87db02bf",
  1496 => x"c288c148",
  1497 => x"d258d4f7",
  1498 => x"d4f7c287",
  1499 => x"87cb02bf",
  1500 => x"bfd0f7c2",
  1501 => x"c280c148",
  1502 => x"c758d4f7",
  1503 => x"d0f7c21e",
  1504 => x"f2c11ebf",
  1505 => x"f6c21ecc",
  1506 => x"49bf97c0",
  1507 => x"497387cc",
  1508 => x"87c8f2c0",
  1509 => x"4b268ef4",
  1510 => x"5e0e4f26",
  1511 => x"0e5d5c5b",
  1512 => x"c086ccff",
  1513 => x"cc59a6e8",
  1514 => x"78c048a6",
  1515 => x"78c080c4",
  1516 => x"78c080c4",
  1517 => x"c8c180c4",
  1518 => x"80c47866",
  1519 => x"80c478c1",
  1520 => x"f7c278c1",
  1521 => x"78c148d4",
  1522 => x"87dfdfff",
  1523 => x"87f8dfff",
  1524 => x"87ccdfff",
  1525 => x"fbc04d70",
  1526 => x"f3c102ad",
  1527 => x"66e4c087",
  1528 => x"87e8c105",
  1529 => x"4a66c4c1",
  1530 => x"7e6a82c4",
  1531 => x"48eccac1",
  1532 => x"4120496e",
  1533 => x"51104120",
  1534 => x"4866c4c1",
  1535 => x"78f2d8c1",
  1536 => x"81c7496a",
  1537 => x"c4c15175",
  1538 => x"81c84966",
  1539 => x"a6dc51c1",
  1540 => x"c178c248",
  1541 => x"c94966c4",
  1542 => x"c151c081",
  1543 => x"ca4966c4",
  1544 => x"c151c081",
  1545 => x"6a1ed81e",
  1546 => x"ff81c849",
  1547 => x"c887edde",
  1548 => x"66c8c186",
  1549 => x"01a8c048",
  1550 => x"a6d487c7",
  1551 => x"cf78c148",
  1552 => x"66c8c187",
  1553 => x"dc88c148",
  1554 => x"87c458a6",
  1555 => x"87f8ddff",
  1556 => x"cb029d75",
  1557 => x"66d487f6",
  1558 => x"66ccc148",
  1559 => x"ebcb03a8",
  1560 => x"ff7ec087",
  1561 => x"7087f9dc",
  1562 => x"c6c1484d",
  1563 => x"58a6c888",
  1564 => x"c1029870",
  1565 => x"c94887d7",
  1566 => x"58a6c888",
  1567 => x"c5029870",
  1568 => x"c14887da",
  1569 => x"58a6c888",
  1570 => x"c2029870",
  1571 => x"c34887f9",
  1572 => x"58a6c888",
  1573 => x"cf029870",
  1574 => x"88c14887",
  1575 => x"7058a6c8",
  1576 => x"f7c40298",
  1577 => x"87c3ca87",
  1578 => x"ff7ef0c0",
  1579 => x"7087f1db",
  1580 => x"adecc04d",
  1581 => x"c487c302",
  1582 => x"ecc05da6",
  1583 => x"87cd02ad",
  1584 => x"87dcdbff",
  1585 => x"ecc04d70",
  1586 => x"f3ff05ad",
  1587 => x"66e4c087",
  1588 => x"87eac105",
  1589 => x"02adecc0",
  1590 => x"dbff87c4",
  1591 => x"1ec087c2",
  1592 => x"66dc1eca",
  1593 => x"c193cc4b",
  1594 => x"c48366cc",
  1595 => x"496c4ca3",
  1596 => x"87e8dbff",
  1597 => x"1ede1ec1",
  1598 => x"dbff496c",
  1599 => x"86d087de",
  1600 => x"7bf2d8c1",
  1601 => x"dc49a3c8",
  1602 => x"a3c95166",
  1603 => x"66e0c049",
  1604 => x"49a3ca51",
  1605 => x"66dc516e",
  1606 => x"c080c148",
  1607 => x"d458a6e0",
  1608 => x"66d84866",
  1609 => x"87cb04a8",
  1610 => x"c14866d4",
  1611 => x"58a6d880",
  1612 => x"d887fec7",
  1613 => x"88c14866",
  1614 => x"c758a6dc",
  1615 => x"daff87f3",
  1616 => x"4d7087c6",
  1617 => x"ff87eac7",
  1618 => x"d087fcdb",
  1619 => x"66d058a6",
  1620 => x"c6c006a8",
  1621 => x"48a6d087",
  1622 => x"ff7866cc",
  1623 => x"c087e8db",
  1624 => x"c105a8ec",
  1625 => x"e4c087f6",
  1626 => x"e6c10566",
  1627 => x"4966d487",
  1628 => x"c4c191cc",
  1629 => x"a1c48166",
  1630 => x"c84c6a4a",
  1631 => x"66cc4aa1",
  1632 => x"ead9c152",
  1633 => x"d7d8ff79",
  1634 => x"9d4d7087",
  1635 => x"c087db02",
  1636 => x"c002adfb",
  1637 => x"547587d4",
  1638 => x"87c4d8ff",
  1639 => x"029d4d70",
  1640 => x"c087c7c0",
  1641 => x"ff05adfb",
  1642 => x"e0c087ec",
  1643 => x"54c1c254",
  1644 => x"d47c97c0",
  1645 => x"66d84866",
  1646 => x"cbc004a8",
  1647 => x"4866d487",
  1648 => x"a6d880c1",
  1649 => x"87e9c558",
  1650 => x"c14866d8",
  1651 => x"58a6dc88",
  1652 => x"ff87dec5",
  1653 => x"7087f1d7",
  1654 => x"87d5c54d",
  1655 => x"c04866cc",
  1656 => x"05a866e4",
  1657 => x"c087f6c4",
  1658 => x"c048a6e8",
  1659 => x"d6d9ff78",
  1660 => x"58a6c487",
  1661 => x"87cfd9ff",
  1662 => x"58a6f0c0",
  1663 => x"05a8ecc0",
  1664 => x"a687c7c0",
  1665 => x"c0786e48",
  1666 => x"d6ff87c4",
  1667 => x"66d487d2",
  1668 => x"c191cc49",
  1669 => x"714866c4",
  1670 => x"58a6c880",
  1671 => x"c84a66c4",
  1672 => x"4966c482",
  1673 => x"516e81ca",
  1674 => x"4966ecc0",
  1675 => x"896e81c1",
  1676 => x"307148c1",
  1677 => x"89c14970",
  1678 => x"c27a9771",
  1679 => x"49bffcf5",
  1680 => x"6a97296e",
  1681 => x"9871484a",
  1682 => x"58a6f4c0",
  1683 => x"c44866c4",
  1684 => x"58a6cc80",
  1685 => x"4cbf66c8",
  1686 => x"4866e4c0",
  1687 => x"02a866cc",
  1688 => x"c087c5c0",
  1689 => x"87c2c07e",
  1690 => x"1e6e7ec1",
  1691 => x"741ee0c0",
  1692 => x"e7d5ff49",
  1693 => x"7086c887",
  1694 => x"adb7c04d",
  1695 => x"87d5c106",
  1696 => x"66c88475",
  1697 => x"e0c049bf",
  1698 => x"4b897481",
  1699 => x"4af8cac1",
  1700 => x"d7defe71",
  1701 => x"c484c287",
  1702 => x"e8c05ca6",
  1703 => x"80c14866",
  1704 => x"58a6ecc0",
  1705 => x"4966f0c0",
  1706 => x"a97081c1",
  1707 => x"87c5c002",
  1708 => x"c2c04cc0",
  1709 => x"744cc187",
  1710 => x"bf66cc1e",
  1711 => x"81e0c049",
  1712 => x"718966c4",
  1713 => x"4966c81e",
  1714 => x"87d0d4ff",
  1715 => x"b7c086c8",
  1716 => x"c5ff01a8",
  1717 => x"66e8c087",
  1718 => x"87d3c002",
  1719 => x"c94966c4",
  1720 => x"66e8c081",
  1721 => x"4866c451",
  1722 => x"78f8dac1",
  1723 => x"c487cec0",
  1724 => x"81c94966",
  1725 => x"66c451c2",
  1726 => x"f6dcc148",
  1727 => x"4866d478",
  1728 => x"04a866d8",
  1729 => x"d487cbc0",
  1730 => x"80c14866",
  1731 => x"c058a6d8",
  1732 => x"66d887d1",
  1733 => x"dc88c148",
  1734 => x"c6c058a6",
  1735 => x"e7d2ff87",
  1736 => x"cc4d7087",
  1737 => x"78c048a6",
  1738 => x"ff87c6c0",
  1739 => x"7087d9d2",
  1740 => x"66e0c04d",
  1741 => x"c080c148",
  1742 => x"7558a6e4",
  1743 => x"cbc0029d",
  1744 => x"4866d487",
  1745 => x"a866ccc1",
  1746 => x"87d5f404",
  1747 => x"c74866d4",
  1748 => x"e1c003a8",
  1749 => x"4c66d487",
  1750 => x"48d4f7c2",
  1751 => x"497478c0",
  1752 => x"c4c191cc",
  1753 => x"a1c48166",
  1754 => x"c04a6a4a",
  1755 => x"84c17952",
  1756 => x"ff04acc7",
  1757 => x"e4c087e2",
  1758 => x"e2c00266",
  1759 => x"66c4c187",
  1760 => x"81d4c149",
  1761 => x"4a66c4c1",
  1762 => x"c082dcc1",
  1763 => x"ead9c152",
  1764 => x"66c4c179",
  1765 => x"81d8c149",
  1766 => x"79fccac1",
  1767 => x"c187d6c0",
  1768 => x"c14966c4",
  1769 => x"c4c181d4",
  1770 => x"d8c14a66",
  1771 => x"c4cbc182",
  1772 => x"e1d9c17a",
  1773 => x"66c4c179",
  1774 => x"81e0c149",
  1775 => x"79c8ddc1",
  1776 => x"87fbcfff",
  1777 => x"ff4866d0",
  1778 => x"4d268ecc",
  1779 => x"4b264c26",
  1780 => x"c71e4f26",
  1781 => x"d0f7c21e",
  1782 => x"f2c11ebf",
  1783 => x"f6c21ecc",
  1784 => x"49bf97c0",
  1785 => x"c187f3ee",
  1786 => x"c049ccf2",
  1787 => x"f487fce1",
  1788 => x"1e4f268e",
  1789 => x"48c0f2c1",
  1790 => x"f3c150c0",
  1791 => x"ff49bff8",
  1792 => x"c087f3d4",
  1793 => x"1e4f2648",
  1794 => x"d4c71e73",
  1795 => x"dcf7c287",
  1796 => x"ff50c048",
  1797 => x"ffc348d4",
  1798 => x"cccbc178",
  1799 => x"f2d6fe49",
  1800 => x"c7e2fe87",
  1801 => x"02987087",
  1802 => x"ebfe87cd",
  1803 => x"987087e5",
  1804 => x"c187c402",
  1805 => x"c087c24a",
  1806 => x"029a724a",
  1807 => x"cbc187c8",
  1808 => x"d6fe49d8",
  1809 => x"f7c287cd",
  1810 => x"78c048d0",
  1811 => x"48c0f6c2",
  1812 => x"fd4950c0",
  1813 => x"dafe87fc",
  1814 => x"9b4b7087",
  1815 => x"c187cf02",
  1816 => x"c75be8f3",
  1817 => x"87f4de49",
  1818 => x"e0c049c1",
  1819 => x"f3c287d0",
  1820 => x"d6e1c087",
  1821 => x"efefc087",
  1822 => x"87f5ff87",
  1823 => x"4f264b26",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000001",
  1827 => x"00001371",
  1828 => x"00002de8",
  1829 => x"44000000",
  1830 => x"00001371",
  1831 => x"00002e06",
  1832 => x"44000000",
  1833 => x"00001371",
  1834 => x"00002e24",
  1835 => x"44000000",
  1836 => x"00001371",
  1837 => x"00002e42",
  1838 => x"44000000",
  1839 => x"00001371",
  1840 => x"00002e60",
  1841 => x"44000000",
  1842 => x"00001371",
  1843 => x"00002e7e",
  1844 => x"44000000",
  1845 => x"00001371",
  1846 => x"00002e9c",
  1847 => x"44000000",
  1848 => x"0000166a",
  1849 => x"00000000",
  1850 => x"44000000",
  1851 => x"00001417",
  1852 => x"00000000",
  1853 => x"44000000",
  1854 => x"000012dc",
  1855 => x"dc86fc1e",
  1856 => x"58a6c487",
  1857 => x"4f268efc",
  1858 => x"48f0fe1e",
  1859 => x"09cd78c0",
  1860 => x"4f260979",
  1861 => x"fcf3c11e",
  1862 => x"2687ed49",
  1863 => x"f0fe1e4f",
  1864 => x"4f2648bf",
  1865 => x"48f0fe1e",
  1866 => x"4f2678c1",
  1867 => x"48f0fe1e",
  1868 => x"4f2678c0",
  1869 => x"c04a711e",
  1870 => x"4f265152",
  1871 => x"5c5b5e0e",
  1872 => x"86f40e5d",
  1873 => x"6d974d71",
  1874 => x"58a6c448",
  1875 => x"974ca5c1",
  1876 => x"a6c8486c",
  1877 => x"c4486e58",
  1878 => x"c505a866",
  1879 => x"c048ff87",
  1880 => x"c7ff87e7",
  1881 => x"49a5c287",
  1882 => x"714b6c97",
  1883 => x"6b974ba3",
  1884 => x"486c974b",
  1885 => x"c158a6c4",
  1886 => x"58a6c880",
  1887 => x"a6cc98c7",
  1888 => x"7c977058",
  1889 => x"7387ddfe",
  1890 => x"268ef448",
  1891 => x"264c264d",
  1892 => x"1e4f264b",
  1893 => x"86f41e73",
  1894 => x"e087d1fe",
  1895 => x"c0494bbf",
  1896 => x"0299c0e0",
  1897 => x"7387ebc0",
  1898 => x"9affc34a",
  1899 => x"97d0fbc2",
  1900 => x"fbc249bf",
  1901 => x"517281d2",
  1902 => x"97d0fbc2",
  1903 => x"a6c448bf",
  1904 => x"c880c158",
  1905 => x"98c758a6",
  1906 => x"c258a6cc",
  1907 => x"c848d0fb",
  1908 => x"c8fd5066",
  1909 => x"58a6c487",
  1910 => x"f487c9fd",
  1911 => x"264b268e",
  1912 => x"fbc21e4f",
  1913 => x"cbfd49d0",
  1914 => x"d3f6c187",
  1915 => x"87d8fc49",
  1916 => x"2687edc4",
  1917 => x"5b5e0e4f",
  1918 => x"fc0e5d5c",
  1919 => x"59a6c486",
  1920 => x"c24dd4ff",
  1921 => x"fc49d0fb",
  1922 => x"4b7087f2",
  1923 => x"04abb7c0",
  1924 => x"c387f8c2",
  1925 => x"c905abf0",
  1926 => x"d8fbc187",
  1927 => x"c278c148",
  1928 => x"e0c387d9",
  1929 => x"87c905ab",
  1930 => x"48dcfbc1",
  1931 => x"cac278c1",
  1932 => x"dcfbc187",
  1933 => x"87c602bf",
  1934 => x"4ca3c0c2",
  1935 => x"4c7387c2",
  1936 => x"bfd8fbc1",
  1937 => x"87e0c002",
  1938 => x"b7c44974",
  1939 => x"fbc19129",
  1940 => x"4a7481e0",
  1941 => x"92c29acf",
  1942 => x"307248c1",
  1943 => x"baff4a70",
  1944 => x"98694872",
  1945 => x"87db7970",
  1946 => x"b7c44974",
  1947 => x"fbc19129",
  1948 => x"4a7481e0",
  1949 => x"92c29acf",
  1950 => x"307248c3",
  1951 => x"69484a70",
  1952 => x"6e7970b0",
  1953 => x"87e7c005",
  1954 => x"c848d0ff",
  1955 => x"7dc578e1",
  1956 => x"bfdcfbc1",
  1957 => x"c387c302",
  1958 => x"fbc17de0",
  1959 => x"c302bfd8",
  1960 => x"7df0c387",
  1961 => x"d0ff7d73",
  1962 => x"78e1c848",
  1963 => x"c178e0c0",
  1964 => x"c048dcfb",
  1965 => x"d8fbc178",
  1966 => x"c278c048",
  1967 => x"f949d0fb",
  1968 => x"4b7087fa",
  1969 => x"03abb7c0",
  1970 => x"c087c8fd",
  1971 => x"268efc48",
  1972 => x"264c264d",
  1973 => x"004f264b",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"54545454",
  1978 => x"54545454",
  1979 => x"54545454",
  1980 => x"54545454",
  1981 => x"54545454",
  1982 => x"54545454",
  1983 => x"54545454",
  1984 => x"54545454",
  1985 => x"54545454",
  1986 => x"54545454",
  1987 => x"54545454",
  1988 => x"54545454",
  1989 => x"54545454",
  1990 => x"54545454",
  1991 => x"54545454",
  1992 => x"724ac01e",
  1993 => x"c191c449",
  1994 => x"c081e0fb",
  1995 => x"d082c179",
  1996 => x"ee04aab7",
  1997 => x"0e4f2687",
  1998 => x"5d5c5b5e",
  1999 => x"f74d710e",
  2000 => x"4a7587ea",
  2001 => x"922ab7c4",
  2002 => x"82e0fbc1",
  2003 => x"9ccf4c75",
  2004 => x"496a94c2",
  2005 => x"c32b744b",
  2006 => x"7448c29b",
  2007 => x"ff4c7030",
  2008 => x"714874bc",
  2009 => x"f67a7098",
  2010 => x"487387fa",
  2011 => x"4c264d26",
  2012 => x"4f264b26",
  2013 => x"48d0ff1e",
  2014 => x"7178e1c8",
  2015 => x"08d4ff48",
  2016 => x"1e4f2678",
  2017 => x"c848d0ff",
  2018 => x"487178e1",
  2019 => x"7808d4ff",
  2020 => x"ff4866c4",
  2021 => x"267808d4",
  2022 => x"4a711e4f",
  2023 => x"1e4966c4",
  2024 => x"deff4972",
  2025 => x"48d0ff87",
  2026 => x"fc78e0c0",
  2027 => x"1e4f268e",
  2028 => x"4b711e73",
  2029 => x"1e4966c8",
  2030 => x"e0c14a73",
  2031 => x"d8ff49a2",
  2032 => x"268efc87",
  2033 => x"1e4f264b",
  2034 => x"c848d0ff",
  2035 => x"487178c9",
  2036 => x"7808d4ff",
  2037 => x"711e4f26",
  2038 => x"87eb494a",
  2039 => x"c848d0ff",
  2040 => x"1e4f2678",
  2041 => x"4b711e73",
  2042 => x"bfe8fbc2",
  2043 => x"c287c302",
  2044 => x"d0ff87eb",
  2045 => x"78c9c848",
  2046 => x"e0c04873",
  2047 => x"08d4ffb0",
  2048 => x"dcfbc278",
  2049 => x"c878c048",
  2050 => x"87c50266",
  2051 => x"c249ffc3",
  2052 => x"c249c087",
  2053 => x"cc59e4fb",
  2054 => x"87c60266",
  2055 => x"4ad5d5c5",
  2056 => x"ffcf87c4",
  2057 => x"fbc24aff",
  2058 => x"fbc25ae8",
  2059 => x"78c148e8",
  2060 => x"4f264b26",
  2061 => x"5c5b5e0e",
  2062 => x"4d710e5d",
  2063 => x"bfe4fbc2",
  2064 => x"029d754b",
  2065 => x"c84987cb",
  2066 => x"dcffc191",
  2067 => x"c482714a",
  2068 => x"dcc3c287",
  2069 => x"124cc04a",
  2070 => x"c2997349",
  2071 => x"48bfe0fb",
  2072 => x"d4ffb871",
  2073 => x"b7c17808",
  2074 => x"b7c8842b",
  2075 => x"87e704ac",
  2076 => x"bfdcfbc2",
  2077 => x"c280c848",
  2078 => x"2658e0fb",
  2079 => x"264c264d",
  2080 => x"1e4f264b",
  2081 => x"4b711e73",
  2082 => x"029a4a13",
  2083 => x"497287cb",
  2084 => x"1387e1fe",
  2085 => x"f5059a4a",
  2086 => x"264b2687",
  2087 => x"fbc21e4f",
  2088 => x"c249bfdc",
  2089 => x"c148dcfb",
  2090 => x"c0c478a1",
  2091 => x"db03a9b7",
  2092 => x"48d4ff87",
  2093 => x"bfe0fbc2",
  2094 => x"dcfbc278",
  2095 => x"fbc249bf",
  2096 => x"a1c148dc",
  2097 => x"b7c0c478",
  2098 => x"87e504a9",
  2099 => x"c848d0ff",
  2100 => x"e8fbc278",
  2101 => x"2678c048",
  2102 => x"0000004f",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"5f000000",
  2106 => x"0000005f",
  2107 => x"00030300",
  2108 => x"00000303",
  2109 => x"147f7f14",
  2110 => x"00147f7f",
  2111 => x"6b2e2400",
  2112 => x"00123a6b",
  2113 => x"18366a4c",
  2114 => x"0032566c",
  2115 => x"594f7e30",
  2116 => x"40683a77",
  2117 => x"07040000",
  2118 => x"00000003",
  2119 => x"3e1c0000",
  2120 => x"00004163",
  2121 => x"63410000",
  2122 => x"00001c3e",
  2123 => x"1c3e2a08",
  2124 => x"082a3e1c",
  2125 => x"3e080800",
  2126 => x"0008083e",
  2127 => x"e0800000",
  2128 => x"00000060",
  2129 => x"08080800",
  2130 => x"00080808",
  2131 => x"60000000",
  2132 => x"00000060",
  2133 => x"18306040",
  2134 => x"0103060c",
  2135 => x"597f3e00",
  2136 => x"003e7f4d",
  2137 => x"7f060400",
  2138 => x"0000007f",
  2139 => x"71634200",
  2140 => x"00464f59",
  2141 => x"49632200",
  2142 => x"00367f49",
  2143 => x"13161c18",
  2144 => x"00107f7f",
  2145 => x"45672700",
  2146 => x"00397d45",
  2147 => x"4b7e3c00",
  2148 => x"00307949",
  2149 => x"71010100",
  2150 => x"00070f79",
  2151 => x"497f3600",
  2152 => x"00367f49",
  2153 => x"494f0600",
  2154 => x"001e3f69",
  2155 => x"66000000",
  2156 => x"00000066",
  2157 => x"e6800000",
  2158 => x"00000066",
  2159 => x"14080800",
  2160 => x"00222214",
  2161 => x"14141400",
  2162 => x"00141414",
  2163 => x"14222200",
  2164 => x"00080814",
  2165 => x"51030200",
  2166 => x"00060f59",
  2167 => x"5d417f3e",
  2168 => x"001e1f55",
  2169 => x"097f7e00",
  2170 => x"007e7f09",
  2171 => x"497f7f00",
  2172 => x"00367f49",
  2173 => x"633e1c00",
  2174 => x"00414141",
  2175 => x"417f7f00",
  2176 => x"001c3e63",
  2177 => x"497f7f00",
  2178 => x"00414149",
  2179 => x"097f7f00",
  2180 => x"00010109",
  2181 => x"417f3e00",
  2182 => x"007a7b49",
  2183 => x"087f7f00",
  2184 => x"007f7f08",
  2185 => x"7f410000",
  2186 => x"0000417f",
  2187 => x"40602000",
  2188 => x"003f7f40",
  2189 => x"1c087f7f",
  2190 => x"00416336",
  2191 => x"407f7f00",
  2192 => x"00404040",
  2193 => x"0c067f7f",
  2194 => x"007f7f06",
  2195 => x"0c067f7f",
  2196 => x"007f7f18",
  2197 => x"417f3e00",
  2198 => x"003e7f41",
  2199 => x"097f7f00",
  2200 => x"00060f09",
  2201 => x"61417f3e",
  2202 => x"00407e7f",
  2203 => x"097f7f00",
  2204 => x"00667f19",
  2205 => x"4d6f2600",
  2206 => x"00327b59",
  2207 => x"7f010100",
  2208 => x"0001017f",
  2209 => x"407f3f00",
  2210 => x"003f7f40",
  2211 => x"703f0f00",
  2212 => x"000f3f70",
  2213 => x"18307f7f",
  2214 => x"007f7f30",
  2215 => x"1c366341",
  2216 => x"4163361c",
  2217 => x"7c060301",
  2218 => x"0103067c",
  2219 => x"4d597161",
  2220 => x"00414347",
  2221 => x"7f7f0000",
  2222 => x"00004141",
  2223 => x"0c060301",
  2224 => x"40603018",
  2225 => x"41410000",
  2226 => x"00007f7f",
  2227 => x"03060c08",
  2228 => x"00080c06",
  2229 => x"80808080",
  2230 => x"00808080",
  2231 => x"03000000",
  2232 => x"00000407",
  2233 => x"54742000",
  2234 => x"00787c54",
  2235 => x"447f7f00",
  2236 => x"00387c44",
  2237 => x"447c3800",
  2238 => x"00004444",
  2239 => x"447c3800",
  2240 => x"007f7f44",
  2241 => x"547c3800",
  2242 => x"00185c54",
  2243 => x"7f7e0400",
  2244 => x"00000505",
  2245 => x"a4bc1800",
  2246 => x"007cfca4",
  2247 => x"047f7f00",
  2248 => x"00787c04",
  2249 => x"3d000000",
  2250 => x"0000407d",
  2251 => x"80808000",
  2252 => x"00007dfd",
  2253 => x"107f7f00",
  2254 => x"00446c38",
  2255 => x"3f000000",
  2256 => x"0000407f",
  2257 => x"180c7c7c",
  2258 => x"00787c0c",
  2259 => x"047c7c00",
  2260 => x"00787c04",
  2261 => x"447c3800",
  2262 => x"00387c44",
  2263 => x"24fcfc00",
  2264 => x"00183c24",
  2265 => x"243c1800",
  2266 => x"00fcfc24",
  2267 => x"047c7c00",
  2268 => x"00080c04",
  2269 => x"545c4800",
  2270 => x"00207454",
  2271 => x"7f3f0400",
  2272 => x"00004444",
  2273 => x"407c3c00",
  2274 => x"007c7c40",
  2275 => x"603c1c00",
  2276 => x"001c3c60",
  2277 => x"30607c3c",
  2278 => x"003c7c60",
  2279 => x"10386c44",
  2280 => x"00446c38",
  2281 => x"e0bc1c00",
  2282 => x"001c3c60",
  2283 => x"74644400",
  2284 => x"00444c5c",
  2285 => x"3e080800",
  2286 => x"00414177",
  2287 => x"7f000000",
  2288 => x"0000007f",
  2289 => x"77414100",
  2290 => x"0008083e",
  2291 => x"03010102",
  2292 => x"00010202",
  2293 => x"7f7f7f7f",
  2294 => x"007f7f7f",
  2295 => x"1c1c0808",
  2296 => x"7f7f3e3e",
  2297 => x"3e3e7f7f",
  2298 => x"08081c1c",
  2299 => x"7c181000",
  2300 => x"0010187c",
  2301 => x"7c301000",
  2302 => x"0010307c",
  2303 => x"60603010",
  2304 => x"00061e78",
  2305 => x"183c6642",
  2306 => x"0042663c",
  2307 => x"c26a3878",
  2308 => x"00386cc6",
  2309 => x"60000060",
  2310 => x"00600000",
  2311 => x"5c5b5e0e",
  2312 => x"86fc0e5d",
  2313 => x"c259a6c4",
  2314 => x"4cbff0fb",
  2315 => x"1ec04bc0",
  2316 => x"02ab66c4",
  2317 => x"4dc087c4",
  2318 => x"4dc187c2",
  2319 => x"49731e75",
  2320 => x"c887e0ee",
  2321 => x"49e0c086",
  2322 => x"c487e9ef",
  2323 => x"496a4aa4",
  2324 => x"f187f0f0",
  2325 => x"84cc87c7",
  2326 => x"b7c883c1",
  2327 => x"cdff04ab",
  2328 => x"268efc87",
  2329 => x"264c264d",
  2330 => x"1e4f264b",
  2331 => x"fbc24a71",
  2332 => x"fbc25af4",
  2333 => x"78c748f4",
  2334 => x"87e0fe49",
  2335 => x"731e4f26",
  2336 => x"fc4b711e",
  2337 => x"730b7b0b",
  2338 => x"c19ac14a",
  2339 => x"ed49a2c0",
  2340 => x"dfc287c4",
  2341 => x"4b265bf4",
  2342 => x"711e4f26",
  2343 => x"1e66c44a",
  2344 => x"caec4972",
  2345 => x"268efc87",
  2346 => x"d4ff1e4f",
  2347 => x"78ffc348",
  2348 => x"c048d0ff",
  2349 => x"d4ff78e1",
  2350 => x"7178c148",
  2351 => x"ff30c448",
  2352 => x"ff7808d4",
  2353 => x"e0c048d0",
  2354 => x"0e4f2678",
  2355 => x"5d5c5b5e",
  2356 => x"c886ec0e",
  2357 => x"78c048a6",
  2358 => x"bfec80c4",
  2359 => x"c280f878",
  2360 => x"78bff0fb",
  2361 => x"bff8fbc2",
  2362 => x"4dbfe84c",
  2363 => x"bff0dfc2",
  2364 => x"87c1e449",
  2365 => x"fee849c7",
  2366 => x"c2497087",
  2367 => x"87d00599",
  2368 => x"bfe8dfc2",
  2369 => x"ccb9ff49",
  2370 => x"99c19966",
  2371 => x"87cdc202",
  2372 => x"ff48a6c8",
  2373 => x"c778bfc8",
  2374 => x"87dbe849",
  2375 => x"a6c44970",
  2376 => x"0599715c",
  2377 => x"66cc87ce",
  2378 => x"c499c149",
  2379 => x"99715ca6",
  2380 => x"87c4c102",
  2381 => x"c84cc8ff",
  2382 => x"a6cc4b66",
  2383 => x"78bfec48",
  2384 => x"cc87f2e2",
  2385 => x"486c5ba6",
  2386 => x"a6d48873",
  2387 => x"a8e8cf58",
  2388 => x"c287d106",
  2389 => x"49bfe4df",
  2390 => x"dfc2b9c1",
  2391 => x"fd7159e8",
  2392 => x"4b6c87c7",
  2393 => x"cee749c7",
  2394 => x"05987087",
  2395 => x"cc87cbff",
  2396 => x"99c14966",
  2397 => x"87c2ff05",
  2398 => x"dfc24c6e",
  2399 => x"c14abff0",
  2400 => x"f4dfc2ba",
  2401 => x"7a0afc5a",
  2402 => x"c19ac10a",
  2403 => x"e949a2c0",
  2404 => x"dac187c4",
  2405 => x"87dfe649",
  2406 => x"c148a6c8",
  2407 => x"e8dfc278",
  2408 => x"7866cc48",
  2409 => x"bff0dfc2",
  2410 => x"87c7c105",
  2411 => x"4bc0c0c8",
  2412 => x"7ed4dfc2",
  2413 => x"49144c6e",
  2414 => x"7087fce5",
  2415 => x"c2c00298",
  2416 => x"c1b57387",
  2417 => x"ff052bb7",
  2418 => x"497587ec",
  2419 => x"7199ffc3",
  2420 => x"fb49c01e",
  2421 => x"497587c4",
  2422 => x"7129b7c8",
  2423 => x"fa49c11e",
  2424 => x"86c887f8",
  2425 => x"e549fdc3",
  2426 => x"fac387cd",
  2427 => x"87c7e549",
  2428 => x"7587d2c7",
  2429 => x"99ffc349",
  2430 => x"712db7c8",
  2431 => x"029d75b5",
  2432 => x"ff87e0c0",
  2433 => x"6e7ebfc8",
  2434 => x"ecdfc249",
  2435 => x"e0c289bf",
  2436 => x"c5c003a9",
  2437 => x"c04dc087",
  2438 => x"dfc287cf",
  2439 => x"786e48ec",
  2440 => x"c287c6c0",
  2441 => x"c048ecdf",
  2442 => x"c8497578",
  2443 => x"cec00599",
  2444 => x"49f5c387",
  2445 => x"7087c0e4",
  2446 => x"0299c249",
  2447 => x"c287ebc0",
  2448 => x"02bff4fb",
  2449 => x"4887cac0",
  2450 => x"fbc288c1",
  2451 => x"d4c058f8",
  2452 => x"4866c487",
  2453 => x"c480e0c1",
  2454 => x"bf6e58a6",
  2455 => x"87c5c002",
  2456 => x"7349ff4b",
  2457 => x"48a6c80f",
  2458 => x"497578c1",
  2459 => x"c00599c4",
  2460 => x"f2c387ce",
  2461 => x"87ffe249",
  2462 => x"99c24970",
  2463 => x"87f2c002",
  2464 => x"bff4fbc2",
  2465 => x"c7486e7e",
  2466 => x"c003a8b7",
  2467 => x"486e87cb",
  2468 => x"fbc280c1",
  2469 => x"d4c058f8",
  2470 => x"4866c487",
  2471 => x"c480e0c1",
  2472 => x"bf6e58a6",
  2473 => x"87c5c002",
  2474 => x"7349fe4b",
  2475 => x"48a6c80f",
  2476 => x"fdc378c1",
  2477 => x"87ffe149",
  2478 => x"99c24970",
  2479 => x"87e6c002",
  2480 => x"bff4fbc2",
  2481 => x"87c9c002",
  2482 => x"48f4fbc2",
  2483 => x"d0c078c0",
  2484 => x"4a66c487",
  2485 => x"6a82e0c1",
  2486 => x"87c5c002",
  2487 => x"7349fd4b",
  2488 => x"48a6c80f",
  2489 => x"fac378c1",
  2490 => x"87cbe149",
  2491 => x"99c24970",
  2492 => x"87eec002",
  2493 => x"bff4fbc2",
  2494 => x"a8b7c748",
  2495 => x"87c9c003",
  2496 => x"48f4fbc2",
  2497 => x"d4c078c7",
  2498 => x"4866c487",
  2499 => x"c480e0c1",
  2500 => x"bf6e58a6",
  2501 => x"87c5c002",
  2502 => x"7349fc4b",
  2503 => x"48a6c80f",
  2504 => x"487578c1",
  2505 => x"c498f0c3",
  2506 => x"987058a6",
  2507 => x"87cec005",
  2508 => x"e049dac1",
  2509 => x"497087c1",
  2510 => x"c10299c2",
  2511 => x"056e87ca",
  2512 => x"c187cdc0",
  2513 => x"dfff49da",
  2514 => x"987087ed",
  2515 => x"87e8c002",
  2516 => x"4b49bfe8",
  2517 => x"c89bffc3",
  2518 => x"b37129b7",
  2519 => x"87d5daff",
  2520 => x"f0c34973",
  2521 => x"05997199",
  2522 => x"c187e5ff",
  2523 => x"dfff49da",
  2524 => x"987087c5",
  2525 => x"87d8ff05",
  2526 => x"bff4fbc2",
  2527 => x"93cc4b49",
  2528 => x"6b8366c4",
  2529 => x"0f73714b",
  2530 => x"c0029c74",
  2531 => x"026c87e9",
  2532 => x"6c87e4c0",
  2533 => x"dedeff49",
  2534 => x"c1497087",
  2535 => x"cbc00299",
  2536 => x"4ba4c487",
  2537 => x"bff4fbc2",
  2538 => x"0f4b6b49",
  2539 => x"c00284c8",
  2540 => x"056c87c5",
  2541 => x"c887dcff",
  2542 => x"c8c00266",
  2543 => x"f4fbc287",
  2544 => x"d7f149bf",
  2545 => x"268eec87",
  2546 => x"264c264d",
  2547 => x"004f264b",
  2548 => x"00000010",
  2549 => x"14111258",
  2550 => x"231c1b1d",
  2551 => x"9491595a",
  2552 => x"f4ebf2f5",
  2553 => x"00000000",
  2554 => x"00000000",
  2555 => x"00000000",
  2556 => x"00000000",
  2557 => x"5c5b5e0e",
  2558 => x"4b710e5d",
  2559 => x"d04cd4ff",
  2560 => x"78c04866",
  2561 => x"ddff49d6",
  2562 => x"ffc387ea",
  2563 => x"c3496c7c",
  2564 => x"4d7199ff",
  2565 => x"99f0c349",
  2566 => x"05a9e0c1",
  2567 => x"ffc387cb",
  2568 => x"c3486c7c",
  2569 => x"0866d098",
  2570 => x"7cffc378",
  2571 => x"c8494a6c",
  2572 => x"7cffc331",
  2573 => x"b2714a6c",
  2574 => x"31c84972",
  2575 => x"6c7cffc3",
  2576 => x"72b2714a",
  2577 => x"c331c849",
  2578 => x"4a6c7cff",
  2579 => x"d0ffb271",
  2580 => x"78e0c048",
  2581 => x"c2029b73",
  2582 => x"757b7287",
  2583 => x"264d2648",
  2584 => x"264b264c",
  2585 => x"4f261e4f",
  2586 => x"5c5b5e0e",
  2587 => x"7686f80e",
  2588 => x"80c4481e",
  2589 => x"fbfd4970",
  2590 => x"7086c487",
  2591 => x"c3486e4b",
  2592 => x"f4c201a8",
  2593 => x"c34a7387",
  2594 => x"d0c19af0",
  2595 => x"87c702aa",
  2596 => x"05aae0c1",
  2597 => x"7387e2c2",
  2598 => x"0299c849",
  2599 => x"c4ff87c3",
  2600 => x"c34c7387",
  2601 => x"05acc29c",
  2602 => x"c487c4c1",
  2603 => x"31c94966",
  2604 => x"66c41e71",
  2605 => x"92ccc14a",
  2606 => x"49fcfbc2",
  2607 => x"ccfe8172",
  2608 => x"49d887fa",
  2609 => x"87ecdaff",
  2610 => x"c21ec0c8",
  2611 => x"fd49f4e8",
  2612 => x"ff87cce6",
  2613 => x"e0c048d0",
  2614 => x"f4e8c278",
  2615 => x"4a66cc1e",
  2616 => x"c292ccc1",
  2617 => x"7249fcfb",
  2618 => x"d0cbfe81",
  2619 => x"c186cc87",
  2620 => x"c4c105ac",
  2621 => x"4966c487",
  2622 => x"1e7131c9",
  2623 => x"c14a66c4",
  2624 => x"fbc292cc",
  2625 => x"817249fc",
  2626 => x"87f0cbfe",
  2627 => x"1ef4e8c2",
  2628 => x"c14a66c8",
  2629 => x"fbc292cc",
  2630 => x"817249fc",
  2631 => x"87dec9fe",
  2632 => x"d9ff49d7",
  2633 => x"c0c887ce",
  2634 => x"f4e8c21e",
  2635 => x"cbe4fd49",
  2636 => x"ff86cc87",
  2637 => x"e0c048d0",
  2638 => x"268ef878",
  2639 => x"264b264c",
  2640 => x"4a711e4f",
  2641 => x"03aab7c4",
  2642 => x"497287ce",
  2643 => x"c291ccc1",
  2644 => x"c181fcfb",
  2645 => x"79c081c8",
  2646 => x"5e0e4f26",
  2647 => x"0e5d5c5b",
  2648 => x"4a7186fc",
  2649 => x"c04bd4ff",
  2650 => x"4d66d44c",
  2651 => x"01adb7c3",
  2652 => x"7287c2c2",
  2653 => x"ecc0029a",
  2654 => x"49751e87",
  2655 => x"c291ccc1",
  2656 => x"7148fcfb",
  2657 => x"58a6c880",
  2658 => x"fe4966c4",
  2659 => x"c487f9c2",
  2660 => x"02987086",
  2661 => x"496e87d4",
  2662 => x"c181c8c1",
  2663 => x"c8496e79",
  2664 => x"c54c6981",
  2665 => x"fe497587",
  2666 => x"d0ff87d7",
  2667 => x"78e1c848",
  2668 => x"48747bdd",
  2669 => x"7098ffc3",
  2670 => x"c849747b",
  2671 => x"487129b7",
  2672 => x"7098ffc3",
  2673 => x"d049747b",
  2674 => x"487129b7",
  2675 => x"7098ffc3",
  2676 => x"d848747b",
  2677 => x"7b7028b7",
  2678 => x"7b7b7bc0",
  2679 => x"7b7b7b7b",
  2680 => x"7b7b7b7b",
  2681 => x"48d0ff7b",
  2682 => x"7578e0c0",
  2683 => x"ff49dc1e",
  2684 => x"c487e6d6",
  2685 => x"268efc86",
  2686 => x"264c264d",
  2687 => x"144f264b",
  2688 => x"1400001d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
