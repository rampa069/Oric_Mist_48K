`define BUILD_DATE "240108"
`define BUILD_TIME "204756"
