
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e4",x"f9",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e4",x"f9",x"c2"),
    14 => (x"48",x"f0",x"e6",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f9",x"e7"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"49",x"72"),
    82 => (x"c2",x"7c",x"71",x"99"),
    83 => (x"05",x"bf",x"f0",x"e6"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"c3",x"29",x"d8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"d0",x"49",x"66",x"d0"),
    90 => (x"99",x"ff",x"c3",x"29"),
    91 => (x"66",x"d0",x"7c",x"71"),
    92 => (x"c3",x"29",x"c8",x"49"),
    93 => (x"7c",x"71",x"99",x"ff"),
    94 => (x"c3",x"49",x"66",x"d0"),
    95 => (x"7c",x"71",x"99",x"ff"),
    96 => (x"29",x"d0",x"49",x"72"),
    97 => (x"71",x"99",x"ff",x"c3"),
    98 => (x"c9",x"4b",x"6c",x"7c"),
    99 => (x"c3",x"4d",x"ff",x"f0"),
   100 => (x"d0",x"05",x"ab",x"ff"),
   101 => (x"7c",x"ff",x"c3",x"87"),
   102 => (x"8d",x"c1",x"4b",x"6c"),
   103 => (x"c3",x"87",x"c6",x"02"),
   104 => (x"f0",x"02",x"ab",x"ff"),
   105 => (x"fe",x"48",x"73",x"87"),
   106 => (x"c0",x"1e",x"87",x"c7"),
   107 => (x"48",x"d4",x"ff",x"49"),
   108 => (x"c1",x"78",x"ff",x"c3"),
   109 => (x"b7",x"c8",x"c3",x"81"),
   110 => (x"87",x"f1",x"04",x"a9"),
   111 => (x"73",x"1e",x"4f",x"26"),
   112 => (x"c4",x"87",x"e7",x"1e"),
   113 => (x"c0",x"4b",x"df",x"f8"),
   114 => (x"f0",x"ff",x"c0",x"1e"),
   115 => (x"fd",x"49",x"f7",x"c1"),
   116 => (x"86",x"c4",x"87",x"e7"),
   117 => (x"c0",x"05",x"a8",x"c1"),
   118 => (x"d4",x"ff",x"87",x"ea"),
   119 => (x"78",x"ff",x"c3",x"48"),
   120 => (x"c0",x"c0",x"c0",x"c1"),
   121 => (x"c0",x"1e",x"c0",x"c0"),
   122 => (x"e9",x"c1",x"f0",x"e1"),
   123 => (x"87",x"c9",x"fd",x"49"),
   124 => (x"98",x"70",x"86",x"c4"),
   125 => (x"ff",x"87",x"ca",x"05"),
   126 => (x"ff",x"c3",x"48",x"d4"),
   127 => (x"cb",x"48",x"c1",x"78"),
   128 => (x"87",x"e6",x"fe",x"87"),
   129 => (x"fe",x"05",x"8b",x"c1"),
   130 => (x"48",x"c0",x"87",x"fd"),
   131 => (x"1e",x"87",x"e6",x"fc"),
   132 => (x"d4",x"ff",x"1e",x"73"),
   133 => (x"78",x"ff",x"c3",x"48"),
   134 => (x"1e",x"c0",x"4b",x"d3"),
   135 => (x"c1",x"f0",x"ff",x"c0"),
   136 => (x"d4",x"fc",x"49",x"c1"),
   137 => (x"70",x"86",x"c4",x"87"),
   138 => (x"87",x"ca",x"05",x"98"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"48",x"c1",x"78",x"ff"),
   141 => (x"f1",x"fd",x"87",x"cb"),
   142 => (x"05",x"8b",x"c1",x"87"),
   143 => (x"c0",x"87",x"db",x"ff"),
   144 => (x"87",x"f1",x"fb",x"48"),
   145 => (x"5c",x"5b",x"5e",x"0e"),
   146 => (x"4c",x"d4",x"ff",x"0e"),
   147 => (x"c6",x"87",x"db",x"fd"),
   148 => (x"e1",x"c0",x"1e",x"ea"),
   149 => (x"49",x"c8",x"c1",x"f0"),
   150 => (x"c4",x"87",x"de",x"fb"),
   151 => (x"02",x"a8",x"c1",x"86"),
   152 => (x"ea",x"fe",x"87",x"c8"),
   153 => (x"c1",x"48",x"c0",x"87"),
   154 => (x"da",x"fa",x"87",x"e2"),
   155 => (x"cf",x"49",x"70",x"87"),
   156 => (x"c6",x"99",x"ff",x"ff"),
   157 => (x"c8",x"02",x"a9",x"ea"),
   158 => (x"87",x"d3",x"fe",x"87"),
   159 => (x"cb",x"c1",x"48",x"c0"),
   160 => (x"7c",x"ff",x"c3",x"87"),
   161 => (x"fc",x"4b",x"f1",x"c0"),
   162 => (x"98",x"70",x"87",x"f4"),
   163 => (x"87",x"eb",x"c0",x"02"),
   164 => (x"ff",x"c0",x"1e",x"c0"),
   165 => (x"49",x"fa",x"c1",x"f0"),
   166 => (x"c4",x"87",x"de",x"fa"),
   167 => (x"05",x"98",x"70",x"86"),
   168 => (x"ff",x"c3",x"87",x"d9"),
   169 => (x"c3",x"49",x"6c",x"7c"),
   170 => (x"7c",x"7c",x"7c",x"ff"),
   171 => (x"99",x"c0",x"c1",x"7c"),
   172 => (x"c1",x"87",x"c4",x"02"),
   173 => (x"c0",x"87",x"d5",x"48"),
   174 => (x"c2",x"87",x"d1",x"48"),
   175 => (x"87",x"c4",x"05",x"ab"),
   176 => (x"87",x"c8",x"48",x"c0"),
   177 => (x"fe",x"05",x"8b",x"c1"),
   178 => (x"48",x"c0",x"87",x"fd"),
   179 => (x"1e",x"87",x"e4",x"f9"),
   180 => (x"e6",x"c2",x"1e",x"73"),
   181 => (x"78",x"c1",x"48",x"f0"),
   182 => (x"d0",x"ff",x"4b",x"c7"),
   183 => (x"fb",x"78",x"c2",x"48"),
   184 => (x"d0",x"ff",x"87",x"c8"),
   185 => (x"c0",x"78",x"c3",x"48"),
   186 => (x"d0",x"e5",x"c0",x"1e"),
   187 => (x"f9",x"49",x"c0",x"c1"),
   188 => (x"86",x"c4",x"87",x"c7"),
   189 => (x"c1",x"05",x"a8",x"c1"),
   190 => (x"ab",x"c2",x"4b",x"87"),
   191 => (x"c0",x"87",x"c5",x"05"),
   192 => (x"87",x"f9",x"c0",x"48"),
   193 => (x"ff",x"05",x"8b",x"c1"),
   194 => (x"f7",x"fc",x"87",x"d0"),
   195 => (x"f4",x"e6",x"c2",x"87"),
   196 => (x"05",x"98",x"70",x"58"),
   197 => (x"1e",x"c1",x"87",x"cd"),
   198 => (x"c1",x"f0",x"ff",x"c0"),
   199 => (x"d8",x"f8",x"49",x"d0"),
   200 => (x"ff",x"86",x"c4",x"87"),
   201 => (x"ff",x"c3",x"48",x"d4"),
   202 => (x"87",x"de",x"c4",x"78"),
   203 => (x"58",x"f8",x"e6",x"c2"),
   204 => (x"c2",x"48",x"d0",x"ff"),
   205 => (x"48",x"d4",x"ff",x"78"),
   206 => (x"c1",x"78",x"ff",x"c3"),
   207 => (x"87",x"f5",x"f7",x"48"),
   208 => (x"5c",x"5b",x"5e",x"0e"),
   209 => (x"4a",x"71",x"0e",x"5d"),
   210 => (x"ff",x"4d",x"ff",x"c3"),
   211 => (x"7c",x"75",x"4c",x"d4"),
   212 => (x"c4",x"48",x"d0",x"ff"),
   213 => (x"7c",x"75",x"78",x"c3"),
   214 => (x"ff",x"c0",x"1e",x"72"),
   215 => (x"49",x"d8",x"c1",x"f0"),
   216 => (x"c4",x"87",x"d6",x"f7"),
   217 => (x"02",x"98",x"70",x"86"),
   218 => (x"48",x"c1",x"87",x"c5"),
   219 => (x"75",x"87",x"f0",x"c0"),
   220 => (x"7c",x"fe",x"c3",x"7c"),
   221 => (x"d4",x"1e",x"c0",x"c8"),
   222 => (x"fa",x"f4",x"49",x"66"),
   223 => (x"75",x"86",x"c4",x"87"),
   224 => (x"75",x"7c",x"75",x"7c"),
   225 => (x"e0",x"da",x"d8",x"7c"),
   226 => (x"6c",x"7c",x"75",x"4b"),
   227 => (x"c5",x"05",x"99",x"49"),
   228 => (x"05",x"8b",x"c1",x"87"),
   229 => (x"7c",x"75",x"87",x"f3"),
   230 => (x"c2",x"48",x"d0",x"ff"),
   231 => (x"f6",x"48",x"c0",x"78"),
   232 => (x"5e",x"0e",x"87",x"cf"),
   233 => (x"0e",x"5d",x"5c",x"5b"),
   234 => (x"4c",x"c0",x"4b",x"71"),
   235 => (x"df",x"cd",x"ee",x"c5"),
   236 => (x"48",x"d4",x"ff",x"4a"),
   237 => (x"68",x"78",x"ff",x"c3"),
   238 => (x"a9",x"fe",x"c3",x"49"),
   239 => (x"87",x"fd",x"c0",x"05"),
   240 => (x"9b",x"73",x"4d",x"70"),
   241 => (x"d0",x"87",x"cc",x"02"),
   242 => (x"49",x"73",x"1e",x"66"),
   243 => (x"c4",x"87",x"cf",x"f4"),
   244 => (x"ff",x"87",x"d6",x"86"),
   245 => (x"d1",x"c4",x"48",x"d0"),
   246 => (x"7d",x"ff",x"c3",x"78"),
   247 => (x"c1",x"48",x"66",x"d0"),
   248 => (x"58",x"a6",x"d4",x"88"),
   249 => (x"f0",x"05",x"98",x"70"),
   250 => (x"48",x"d4",x"ff",x"87"),
   251 => (x"78",x"78",x"ff",x"c3"),
   252 => (x"c5",x"05",x"9b",x"73"),
   253 => (x"48",x"d0",x"ff",x"87"),
   254 => (x"4a",x"c1",x"78",x"d0"),
   255 => (x"05",x"8a",x"c1",x"4c"),
   256 => (x"74",x"87",x"ee",x"fe"),
   257 => (x"87",x"e9",x"f4",x"48"),
   258 => (x"71",x"1e",x"73",x"1e"),
   259 => (x"ff",x"4b",x"c0",x"4a"),
   260 => (x"ff",x"c3",x"48",x"d4"),
   261 => (x"48",x"d0",x"ff",x"78"),
   262 => (x"ff",x"78",x"c3",x"c4"),
   263 => (x"ff",x"c3",x"48",x"d4"),
   264 => (x"c0",x"1e",x"72",x"78"),
   265 => (x"d1",x"c1",x"f0",x"ff"),
   266 => (x"87",x"cd",x"f4",x"49"),
   267 => (x"98",x"70",x"86",x"c4"),
   268 => (x"c8",x"87",x"d2",x"05"),
   269 => (x"66",x"cc",x"1e",x"c0"),
   270 => (x"87",x"e6",x"fd",x"49"),
   271 => (x"4b",x"70",x"86",x"c4"),
   272 => (x"c2",x"48",x"d0",x"ff"),
   273 => (x"f3",x"48",x"73",x"78"),
   274 => (x"5e",x"0e",x"87",x"eb"),
   275 => (x"0e",x"5d",x"5c",x"5b"),
   276 => (x"ff",x"c0",x"1e",x"c0"),
   277 => (x"49",x"c9",x"c1",x"f0"),
   278 => (x"d2",x"87",x"de",x"f3"),
   279 => (x"f8",x"e6",x"c2",x"1e"),
   280 => (x"87",x"fe",x"fc",x"49"),
   281 => (x"4c",x"c0",x"86",x"c8"),
   282 => (x"b7",x"d2",x"84",x"c1"),
   283 => (x"87",x"f8",x"04",x"ac"),
   284 => (x"97",x"f8",x"e6",x"c2"),
   285 => (x"c0",x"c3",x"49",x"bf"),
   286 => (x"a9",x"c0",x"c1",x"99"),
   287 => (x"87",x"e7",x"c0",x"05"),
   288 => (x"97",x"ff",x"e6",x"c2"),
   289 => (x"31",x"d0",x"49",x"bf"),
   290 => (x"97",x"c0",x"e7",x"c2"),
   291 => (x"32",x"c8",x"4a",x"bf"),
   292 => (x"e7",x"c2",x"b1",x"72"),
   293 => (x"4a",x"bf",x"97",x"c1"),
   294 => (x"cf",x"4c",x"71",x"b1"),
   295 => (x"9c",x"ff",x"ff",x"ff"),
   296 => (x"34",x"ca",x"84",x"c1"),
   297 => (x"c2",x"87",x"e7",x"c1"),
   298 => (x"bf",x"97",x"c1",x"e7"),
   299 => (x"c6",x"31",x"c1",x"49"),
   300 => (x"c2",x"e7",x"c2",x"99"),
   301 => (x"c7",x"4a",x"bf",x"97"),
   302 => (x"b1",x"72",x"2a",x"b7"),
   303 => (x"97",x"fd",x"e6",x"c2"),
   304 => (x"cf",x"4d",x"4a",x"bf"),
   305 => (x"fe",x"e6",x"c2",x"9d"),
   306 => (x"c3",x"4a",x"bf",x"97"),
   307 => (x"c2",x"32",x"ca",x"9a"),
   308 => (x"bf",x"97",x"ff",x"e6"),
   309 => (x"73",x"33",x"c2",x"4b"),
   310 => (x"c0",x"e7",x"c2",x"b2"),
   311 => (x"c3",x"4b",x"bf",x"97"),
   312 => (x"b7",x"c6",x"9b",x"c0"),
   313 => (x"c2",x"b2",x"73",x"2b"),
   314 => (x"71",x"48",x"c1",x"81"),
   315 => (x"c1",x"49",x"70",x"30"),
   316 => (x"70",x"30",x"75",x"48"),
   317 => (x"c1",x"4c",x"72",x"4d"),
   318 => (x"c8",x"94",x"71",x"84"),
   319 => (x"06",x"ad",x"b7",x"c0"),
   320 => (x"34",x"c1",x"87",x"cc"),
   321 => (x"c0",x"c8",x"2d",x"b7"),
   322 => (x"ff",x"01",x"ad",x"b7"),
   323 => (x"48",x"74",x"87",x"f4"),
   324 => (x"0e",x"87",x"de",x"f0"),
   325 => (x"5d",x"5c",x"5b",x"5e"),
   326 => (x"c2",x"86",x"f8",x"0e"),
   327 => (x"c0",x"48",x"de",x"ef"),
   328 => (x"d6",x"e7",x"c2",x"78"),
   329 => (x"fb",x"49",x"c0",x"1e"),
   330 => (x"86",x"c4",x"87",x"de"),
   331 => (x"c5",x"05",x"98",x"70"),
   332 => (x"c9",x"48",x"c0",x"87"),
   333 => (x"4d",x"c0",x"87",x"ce"),
   334 => (x"f2",x"c0",x"7e",x"c1"),
   335 => (x"c2",x"49",x"bf",x"ed"),
   336 => (x"71",x"4a",x"cc",x"e8"),
   337 => (x"e0",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"7e",x"c0",x"87",x"c2"),
   340 => (x"bf",x"e9",x"f2",x"c0"),
   341 => (x"e8",x"e8",x"c2",x"49"),
   342 => (x"4b",x"c8",x"71",x"4a"),
   343 => (x"70",x"87",x"ca",x"ec"),
   344 => (x"87",x"c2",x"05",x"98"),
   345 => (x"02",x"6e",x"7e",x"c0"),
   346 => (x"c2",x"87",x"fd",x"c0"),
   347 => (x"4d",x"bf",x"dc",x"ee"),
   348 => (x"9f",x"d4",x"ef",x"c2"),
   349 => (x"c5",x"48",x"7e",x"bf"),
   350 => (x"05",x"a8",x"ea",x"d6"),
   351 => (x"ee",x"c2",x"87",x"c7"),
   352 => (x"ce",x"4d",x"bf",x"dc"),
   353 => (x"ca",x"48",x"6e",x"87"),
   354 => (x"02",x"a8",x"d5",x"e9"),
   355 => (x"48",x"c0",x"87",x"c5"),
   356 => (x"c2",x"87",x"f1",x"c7"),
   357 => (x"75",x"1e",x"d6",x"e7"),
   358 => (x"87",x"ec",x"f9",x"49"),
   359 => (x"98",x"70",x"86",x"c4"),
   360 => (x"c0",x"87",x"c5",x"05"),
   361 => (x"87",x"dc",x"c7",x"48"),
   362 => (x"bf",x"e9",x"f2",x"c0"),
   363 => (x"e8",x"e8",x"c2",x"49"),
   364 => (x"4b",x"c8",x"71",x"4a"),
   365 => (x"70",x"87",x"f2",x"ea"),
   366 => (x"87",x"c8",x"05",x"98"),
   367 => (x"48",x"de",x"ef",x"c2"),
   368 => (x"87",x"da",x"78",x"c1"),
   369 => (x"bf",x"ed",x"f2",x"c0"),
   370 => (x"cc",x"e8",x"c2",x"49"),
   371 => (x"4b",x"c8",x"71",x"4a"),
   372 => (x"70",x"87",x"d6",x"ea"),
   373 => (x"c5",x"c0",x"02",x"98"),
   374 => (x"c6",x"48",x"c0",x"87"),
   375 => (x"ef",x"c2",x"87",x"e6"),
   376 => (x"49",x"bf",x"97",x"d4"),
   377 => (x"05",x"a9",x"d5",x"c1"),
   378 => (x"c2",x"87",x"cd",x"c0"),
   379 => (x"bf",x"97",x"d5",x"ef"),
   380 => (x"a9",x"ea",x"c2",x"49"),
   381 => (x"87",x"c5",x"c0",x"02"),
   382 => (x"c7",x"c6",x"48",x"c0"),
   383 => (x"d6",x"e7",x"c2",x"87"),
   384 => (x"48",x"7e",x"bf",x"97"),
   385 => (x"02",x"a8",x"e9",x"c3"),
   386 => (x"6e",x"87",x"ce",x"c0"),
   387 => (x"a8",x"eb",x"c3",x"48"),
   388 => (x"87",x"c5",x"c0",x"02"),
   389 => (x"eb",x"c5",x"48",x"c0"),
   390 => (x"e1",x"e7",x"c2",x"87"),
   391 => (x"99",x"49",x"bf",x"97"),
   392 => (x"87",x"cc",x"c0",x"05"),
   393 => (x"97",x"e2",x"e7",x"c2"),
   394 => (x"a9",x"c2",x"49",x"bf"),
   395 => (x"87",x"c5",x"c0",x"02"),
   396 => (x"cf",x"c5",x"48",x"c0"),
   397 => (x"e3",x"e7",x"c2",x"87"),
   398 => (x"c2",x"48",x"bf",x"97"),
   399 => (x"70",x"58",x"da",x"ef"),
   400 => (x"88",x"c1",x"48",x"4c"),
   401 => (x"58",x"de",x"ef",x"c2"),
   402 => (x"97",x"e4",x"e7",x"c2"),
   403 => (x"81",x"75",x"49",x"bf"),
   404 => (x"97",x"e5",x"e7",x"c2"),
   405 => (x"32",x"c8",x"4a",x"bf"),
   406 => (x"c2",x"7e",x"a1",x"72"),
   407 => (x"6e",x"48",x"eb",x"f3"),
   408 => (x"e6",x"e7",x"c2",x"78"),
   409 => (x"c8",x"48",x"bf",x"97"),
   410 => (x"ef",x"c2",x"58",x"a6"),
   411 => (x"c2",x"02",x"bf",x"de"),
   412 => (x"f2",x"c0",x"87",x"d4"),
   413 => (x"c2",x"49",x"bf",x"e9"),
   414 => (x"71",x"4a",x"e8",x"e8"),
   415 => (x"e8",x"e7",x"4b",x"c8"),
   416 => (x"02",x"98",x"70",x"87"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"f8",x"c3",x"48"),
   419 => (x"bf",x"d6",x"ef",x"c2"),
   420 => (x"ff",x"f3",x"c2",x"4c"),
   421 => (x"fb",x"e7",x"c2",x"5c"),
   422 => (x"c8",x"49",x"bf",x"97"),
   423 => (x"fa",x"e7",x"c2",x"31"),
   424 => (x"a1",x"4a",x"bf",x"97"),
   425 => (x"fc",x"e7",x"c2",x"49"),
   426 => (x"d0",x"4a",x"bf",x"97"),
   427 => (x"49",x"a1",x"72",x"32"),
   428 => (x"97",x"fd",x"e7",x"c2"),
   429 => (x"32",x"d8",x"4a",x"bf"),
   430 => (x"c4",x"49",x"a1",x"72"),
   431 => (x"f3",x"c2",x"91",x"66"),
   432 => (x"c2",x"81",x"bf",x"eb"),
   433 => (x"c2",x"59",x"f3",x"f3"),
   434 => (x"bf",x"97",x"c3",x"e8"),
   435 => (x"c2",x"32",x"c8",x"4a"),
   436 => (x"bf",x"97",x"c2",x"e8"),
   437 => (x"c2",x"4a",x"a2",x"4b"),
   438 => (x"bf",x"97",x"c4",x"e8"),
   439 => (x"73",x"33",x"d0",x"4b"),
   440 => (x"e8",x"c2",x"4a",x"a2"),
   441 => (x"4b",x"bf",x"97",x"c5"),
   442 => (x"33",x"d8",x"9b",x"cf"),
   443 => (x"c2",x"4a",x"a2",x"73"),
   444 => (x"c2",x"5a",x"f7",x"f3"),
   445 => (x"4a",x"bf",x"f3",x"f3"),
   446 => (x"92",x"74",x"8a",x"c2"),
   447 => (x"48",x"f7",x"f3",x"c2"),
   448 => (x"c1",x"78",x"a1",x"72"),
   449 => (x"e7",x"c2",x"87",x"ca"),
   450 => (x"49",x"bf",x"97",x"e8"),
   451 => (x"e7",x"c2",x"31",x"c8"),
   452 => (x"4a",x"bf",x"97",x"e7"),
   453 => (x"ef",x"c2",x"49",x"a1"),
   454 => (x"ef",x"c2",x"59",x"e6"),
   455 => (x"c5",x"49",x"bf",x"e2"),
   456 => (x"81",x"ff",x"c7",x"31"),
   457 => (x"f3",x"c2",x"29",x"c9"),
   458 => (x"e7",x"c2",x"59",x"ff"),
   459 => (x"4a",x"bf",x"97",x"ed"),
   460 => (x"e7",x"c2",x"32",x"c8"),
   461 => (x"4b",x"bf",x"97",x"ec"),
   462 => (x"66",x"c4",x"4a",x"a2"),
   463 => (x"c2",x"82",x"6e",x"92"),
   464 => (x"c2",x"5a",x"fb",x"f3"),
   465 => (x"c0",x"48",x"f3",x"f3"),
   466 => (x"ef",x"f3",x"c2",x"78"),
   467 => (x"78",x"a1",x"72",x"48"),
   468 => (x"48",x"ff",x"f3",x"c2"),
   469 => (x"bf",x"f3",x"f3",x"c2"),
   470 => (x"c3",x"f4",x"c2",x"78"),
   471 => (x"f7",x"f3",x"c2",x"48"),
   472 => (x"ef",x"c2",x"78",x"bf"),
   473 => (x"c0",x"02",x"bf",x"de"),
   474 => (x"48",x"74",x"87",x"c9"),
   475 => (x"7e",x"70",x"30",x"c4"),
   476 => (x"c2",x"87",x"c9",x"c0"),
   477 => (x"48",x"bf",x"fb",x"f3"),
   478 => (x"7e",x"70",x"30",x"c4"),
   479 => (x"48",x"e2",x"ef",x"c2"),
   480 => (x"48",x"c1",x"78",x"6e"),
   481 => (x"4d",x"26",x"8e",x"f8"),
   482 => (x"4b",x"26",x"4c",x"26"),
   483 => (x"5e",x"0e",x"4f",x"26"),
   484 => (x"0e",x"5d",x"5c",x"5b"),
   485 => (x"ef",x"c2",x"4a",x"71"),
   486 => (x"cb",x"02",x"bf",x"de"),
   487 => (x"c7",x"4b",x"72",x"87"),
   488 => (x"c1",x"4c",x"72",x"2b"),
   489 => (x"87",x"c9",x"9c",x"ff"),
   490 => (x"2b",x"c8",x"4b",x"72"),
   491 => (x"ff",x"c3",x"4c",x"72"),
   492 => (x"eb",x"f3",x"c2",x"9c"),
   493 => (x"f2",x"c0",x"83",x"bf"),
   494 => (x"02",x"ab",x"bf",x"e5"),
   495 => (x"f2",x"c0",x"87",x"d9"),
   496 => (x"e7",x"c2",x"5b",x"e9"),
   497 => (x"49",x"73",x"1e",x"d6"),
   498 => (x"c4",x"87",x"fd",x"f0"),
   499 => (x"05",x"98",x"70",x"86"),
   500 => (x"48",x"c0",x"87",x"c5"),
   501 => (x"c2",x"87",x"e6",x"c0"),
   502 => (x"02",x"bf",x"de",x"ef"),
   503 => (x"49",x"74",x"87",x"d2"),
   504 => (x"e7",x"c2",x"91",x"c4"),
   505 => (x"4d",x"69",x"81",x"d6"),
   506 => (x"ff",x"ff",x"ff",x"cf"),
   507 => (x"87",x"cb",x"9d",x"ff"),
   508 => (x"91",x"c2",x"49",x"74"),
   509 => (x"81",x"d6",x"e7",x"c2"),
   510 => (x"75",x"4d",x"69",x"9f"),
   511 => (x"87",x"c6",x"fe",x"48"),
   512 => (x"5c",x"5b",x"5e",x"0e"),
   513 => (x"86",x"f8",x"0e",x"5d"),
   514 => (x"05",x"9c",x"4c",x"71"),
   515 => (x"48",x"c0",x"87",x"c5"),
   516 => (x"c8",x"87",x"c2",x"c3"),
   517 => (x"48",x"6e",x"7e",x"a4"),
   518 => (x"66",x"d8",x"78",x"c0"),
   519 => (x"d8",x"87",x"c7",x"02"),
   520 => (x"05",x"bf",x"97",x"66"),
   521 => (x"48",x"c0",x"87",x"c5"),
   522 => (x"c0",x"87",x"ea",x"c2"),
   523 => (x"49",x"49",x"c1",x"1e"),
   524 => (x"c4",x"87",x"d7",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"e6",x"ef",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c8"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ed"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"d5",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"de",x"ef"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ec"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"da",x"ef",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fb",x"f9"),
   581 => (x"d6",x"ef",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"da",x"ef",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d2",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"ef",x"f3",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"d6",x"ef",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"da",x"ef",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"e9",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d5",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c7",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"ef",x"f3",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"d6",x"ef",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"da",x"ef",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"e9"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"fe"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f8"),
   629 => (x"0e",x"5d",x"5c",x"5b"),
   630 => (x"d4",x"4b",x"71",x"1e"),
   631 => (x"9b",x"73",x"4d",x"66"),
   632 => (x"87",x"cc",x"c1",x"02"),
   633 => (x"69",x"49",x"a3",x"c8"),
   634 => (x"87",x"c4",x"c1",x"02"),
   635 => (x"c2",x"4c",x"a3",x"d0"),
   636 => (x"49",x"bf",x"da",x"ef"),
   637 => (x"4a",x"6c",x"b9",x"ff"),
   638 => (x"66",x"d4",x"7e",x"99"),
   639 => (x"87",x"cd",x"06",x"a9"),
   640 => (x"cc",x"7c",x"7b",x"c0"),
   641 => (x"a3",x"c4",x"4a",x"a3"),
   642 => (x"ca",x"79",x"6a",x"49"),
   643 => (x"f8",x"49",x"72",x"87"),
   644 => (x"66",x"d4",x"99",x"c0"),
   645 => (x"75",x"8d",x"71",x"4d"),
   646 => (x"71",x"29",x"c9",x"49"),
   647 => (x"fa",x"49",x"73",x"1e"),
   648 => (x"e7",x"c2",x"87",x"f8"),
   649 => (x"49",x"73",x"1e",x"d6"),
   650 => (x"c8",x"87",x"c9",x"fc"),
   651 => (x"7c",x"66",x"d4",x"86"),
   652 => (x"87",x"d2",x"f5",x"26"),
   653 => (x"71",x"1e",x"73",x"1e"),
   654 => (x"c0",x"02",x"9b",x"4b"),
   655 => (x"f4",x"c2",x"87",x"e4"),
   656 => (x"4a",x"73",x"5b",x"c3"),
   657 => (x"ef",x"c2",x"8a",x"c2"),
   658 => (x"92",x"49",x"bf",x"d6"),
   659 => (x"bf",x"ef",x"f3",x"c2"),
   660 => (x"c2",x"80",x"72",x"48"),
   661 => (x"71",x"58",x"c7",x"f4"),
   662 => (x"c2",x"30",x"c4",x"48"),
   663 => (x"c0",x"58",x"e6",x"ef"),
   664 => (x"f3",x"c2",x"87",x"ed"),
   665 => (x"f3",x"c2",x"48",x"ff"),
   666 => (x"c2",x"78",x"bf",x"f3"),
   667 => (x"c2",x"48",x"c3",x"f4"),
   668 => (x"78",x"bf",x"f7",x"f3"),
   669 => (x"bf",x"de",x"ef",x"c2"),
   670 => (x"c2",x"87",x"c9",x"02"),
   671 => (x"49",x"bf",x"d6",x"ef"),
   672 => (x"87",x"c7",x"31",x"c4"),
   673 => (x"bf",x"fb",x"f3",x"c2"),
   674 => (x"c2",x"31",x"c4",x"49"),
   675 => (x"f3",x"59",x"e6",x"ef"),
   676 => (x"5e",x"0e",x"87",x"f8"),
   677 => (x"71",x"0e",x"5c",x"5b"),
   678 => (x"72",x"4b",x"c0",x"4a"),
   679 => (x"e1",x"c0",x"02",x"9a"),
   680 => (x"49",x"a2",x"da",x"87"),
   681 => (x"c2",x"4b",x"69",x"9f"),
   682 => (x"02",x"bf",x"de",x"ef"),
   683 => (x"a2",x"d4",x"87",x"cf"),
   684 => (x"49",x"69",x"9f",x"49"),
   685 => (x"ff",x"ff",x"c0",x"4c"),
   686 => (x"c2",x"34",x"d0",x"9c"),
   687 => (x"74",x"4c",x"c0",x"87"),
   688 => (x"49",x"73",x"b3",x"49"),
   689 => (x"f2",x"87",x"ed",x"fd"),
   690 => (x"5e",x"0e",x"87",x"fe"),
   691 => (x"0e",x"5d",x"5c",x"5b"),
   692 => (x"4a",x"71",x"86",x"f4"),
   693 => (x"9a",x"72",x"7e",x"c0"),
   694 => (x"c2",x"87",x"d8",x"02"),
   695 => (x"c0",x"48",x"d2",x"e7"),
   696 => (x"ca",x"e7",x"c2",x"78"),
   697 => (x"c3",x"f4",x"c2",x"48"),
   698 => (x"e7",x"c2",x"78",x"bf"),
   699 => (x"f3",x"c2",x"48",x"ce"),
   700 => (x"c2",x"78",x"bf",x"ff"),
   701 => (x"c0",x"48",x"f3",x"ef"),
   702 => (x"e2",x"ef",x"c2",x"50"),
   703 => (x"e7",x"c2",x"49",x"bf"),
   704 => (x"71",x"4a",x"bf",x"d2"),
   705 => (x"c9",x"c4",x"03",x"aa"),
   706 => (x"cf",x"49",x"72",x"87"),
   707 => (x"e9",x"c0",x"05",x"99"),
   708 => (x"e5",x"f2",x"c0",x"87"),
   709 => (x"ca",x"e7",x"c2",x"48"),
   710 => (x"e7",x"c2",x"78",x"bf"),
   711 => (x"e7",x"c2",x"1e",x"d6"),
   712 => (x"c2",x"49",x"bf",x"ca"),
   713 => (x"c1",x"48",x"ca",x"e7"),
   714 => (x"e3",x"71",x"78",x"a1"),
   715 => (x"86",x"c4",x"87",x"da"),
   716 => (x"48",x"e1",x"f2",x"c0"),
   717 => (x"78",x"d6",x"e7",x"c2"),
   718 => (x"f2",x"c0",x"87",x"cc"),
   719 => (x"c0",x"48",x"bf",x"e1"),
   720 => (x"f2",x"c0",x"80",x"e0"),
   721 => (x"e7",x"c2",x"58",x"e5"),
   722 => (x"c1",x"48",x"bf",x"d2"),
   723 => (x"d6",x"e7",x"c2",x"80"),
   724 => (x"0c",x"a1",x"27",x"58"),
   725 => (x"97",x"bf",x"00",x"00"),
   726 => (x"02",x"9d",x"4d",x"bf"),
   727 => (x"c3",x"87",x"e3",x"c2"),
   728 => (x"c2",x"02",x"ad",x"e5"),
   729 => (x"f2",x"c0",x"87",x"dc"),
   730 => (x"cb",x"4b",x"bf",x"e1"),
   731 => (x"4c",x"11",x"49",x"a3"),
   732 => (x"c1",x"05",x"ac",x"cf"),
   733 => (x"49",x"75",x"87",x"d2"),
   734 => (x"89",x"c1",x"99",x"df"),
   735 => (x"ef",x"c2",x"91",x"cd"),
   736 => (x"a3",x"c1",x"81",x"e6"),
   737 => (x"c3",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"c5"),
   740 => (x"4a",x"a3",x"c7",x"51"),
   741 => (x"a3",x"c9",x"51",x"12"),
   742 => (x"ce",x"51",x"12",x"4a"),
   743 => (x"51",x"12",x"4a",x"a3"),
   744 => (x"12",x"4a",x"a3",x"d0"),
   745 => (x"4a",x"a3",x"d2",x"51"),
   746 => (x"a3",x"d4",x"51",x"12"),
   747 => (x"d6",x"51",x"12",x"4a"),
   748 => (x"51",x"12",x"4a",x"a3"),
   749 => (x"12",x"4a",x"a3",x"d8"),
   750 => (x"4a",x"a3",x"dc",x"51"),
   751 => (x"a3",x"de",x"51",x"12"),
   752 => (x"c1",x"51",x"12",x"4a"),
   753 => (x"87",x"fa",x"c0",x"7e"),
   754 => (x"99",x"c8",x"49",x"74"),
   755 => (x"87",x"eb",x"c0",x"05"),
   756 => (x"99",x"d0",x"49",x"74"),
   757 => (x"dc",x"87",x"d1",x"05"),
   758 => (x"cb",x"c0",x"02",x"66"),
   759 => (x"dc",x"49",x"73",x"87"),
   760 => (x"98",x"70",x"0f",x"66"),
   761 => (x"87",x"d3",x"c0",x"02"),
   762 => (x"c6",x"c0",x"05",x"6e"),
   763 => (x"e6",x"ef",x"c2",x"87"),
   764 => (x"c0",x"50",x"c0",x"48"),
   765 => (x"48",x"bf",x"e1",x"f2"),
   766 => (x"c2",x"87",x"e1",x"c2"),
   767 => (x"c0",x"48",x"f3",x"ef"),
   768 => (x"ef",x"c2",x"7e",x"50"),
   769 => (x"c2",x"49",x"bf",x"e2"),
   770 => (x"4a",x"bf",x"d2",x"e7"),
   771 => (x"fb",x"04",x"aa",x"71"),
   772 => (x"f4",x"c2",x"87",x"f7"),
   773 => (x"c0",x"05",x"bf",x"c3"),
   774 => (x"ef",x"c2",x"87",x"c8"),
   775 => (x"c1",x"02",x"bf",x"de"),
   776 => (x"e7",x"c2",x"87",x"f8"),
   777 => (x"ed",x"49",x"bf",x"ce"),
   778 => (x"49",x"70",x"87",x"e4"),
   779 => (x"59",x"d2",x"e7",x"c2"),
   780 => (x"c2",x"48",x"a6",x"c4"),
   781 => (x"78",x"bf",x"ce",x"e7"),
   782 => (x"bf",x"de",x"ef",x"c2"),
   783 => (x"87",x"d8",x"c0",x"02"),
   784 => (x"cf",x"49",x"66",x"c4"),
   785 => (x"f8",x"ff",x"ff",x"ff"),
   786 => (x"c0",x"02",x"a9",x"99"),
   787 => (x"4c",x"c0",x"87",x"c5"),
   788 => (x"c1",x"87",x"e1",x"c0"),
   789 => (x"87",x"dc",x"c0",x"4c"),
   790 => (x"cf",x"49",x"66",x"c4"),
   791 => (x"a9",x"99",x"f8",x"ff"),
   792 => (x"87",x"c8",x"c0",x"02"),
   793 => (x"c0",x"48",x"a6",x"c8"),
   794 => (x"87",x"c5",x"c0",x"78"),
   795 => (x"c1",x"48",x"a6",x"c8"),
   796 => (x"4c",x"66",x"c8",x"78"),
   797 => (x"c0",x"05",x"9c",x"74"),
   798 => (x"66",x"c4",x"87",x"e0"),
   799 => (x"c2",x"89",x"c2",x"49"),
   800 => (x"4a",x"bf",x"d6",x"ef"),
   801 => (x"ef",x"f3",x"c2",x"91"),
   802 => (x"e7",x"c2",x"4a",x"bf"),
   803 => (x"a1",x"72",x"48",x"ca"),
   804 => (x"d2",x"e7",x"c2",x"78"),
   805 => (x"f9",x"78",x"c0",x"48"),
   806 => (x"48",x"c0",x"87",x"df"),
   807 => (x"e5",x"eb",x"8e",x"f4"),
   808 => (x"00",x"00",x"00",x"87"),
   809 => (x"ff",x"ff",x"ff",x"00"),
   810 => (x"00",x"0c",x"b1",x"ff"),
   811 => (x"00",x"0c",x"ba",x"00"),
   812 => (x"54",x"41",x"46",x"00"),
   813 => (x"20",x"20",x"32",x"33"),
   814 => (x"41",x"46",x"00",x"20"),
   815 => (x"20",x"36",x"31",x"54"),
   816 => (x"1e",x"00",x"20",x"20"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"48",x"68",x"78",x"ff"),
   819 => (x"ff",x"1e",x"4f",x"26"),
   820 => (x"ff",x"c3",x"48",x"d4"),
   821 => (x"48",x"d0",x"ff",x"78"),
   822 => (x"ff",x"78",x"e1",x"c0"),
   823 => (x"78",x"d4",x"48",x"d4"),
   824 => (x"48",x"c7",x"f4",x"c2"),
   825 => (x"50",x"bf",x"d4",x"ff"),
   826 => (x"ff",x"1e",x"4f",x"26"),
   827 => (x"e0",x"c0",x"48",x"d0"),
   828 => (x"1e",x"4f",x"26",x"78"),
   829 => (x"70",x"87",x"cc",x"ff"),
   830 => (x"c6",x"02",x"99",x"49"),
   831 => (x"a9",x"fb",x"c0",x"87"),
   832 => (x"71",x"87",x"f1",x"05"),
   833 => (x"0e",x"4f",x"26",x"48"),
   834 => (x"0e",x"5c",x"5b",x"5e"),
   835 => (x"4c",x"c0",x"4b",x"71"),
   836 => (x"70",x"87",x"f0",x"fe"),
   837 => (x"c0",x"02",x"99",x"49"),
   838 => (x"ec",x"c0",x"87",x"f9"),
   839 => (x"f2",x"c0",x"02",x"a9"),
   840 => (x"a9",x"fb",x"c0",x"87"),
   841 => (x"87",x"eb",x"c0",x"02"),
   842 => (x"ac",x"b7",x"66",x"cc"),
   843 => (x"d0",x"87",x"c7",x"03"),
   844 => (x"87",x"c2",x"02",x"66"),
   845 => (x"99",x"71",x"53",x"71"),
   846 => (x"c1",x"87",x"c2",x"02"),
   847 => (x"87",x"c3",x"fe",x"84"),
   848 => (x"02",x"99",x"49",x"70"),
   849 => (x"ec",x"c0",x"87",x"cd"),
   850 => (x"87",x"c7",x"02",x"a9"),
   851 => (x"05",x"a9",x"fb",x"c0"),
   852 => (x"d0",x"87",x"d5",x"ff"),
   853 => (x"87",x"c3",x"02",x"66"),
   854 => (x"c0",x"7b",x"97",x"c0"),
   855 => (x"c4",x"05",x"a9",x"ec"),
   856 => (x"c5",x"4a",x"74",x"87"),
   857 => (x"c0",x"4a",x"74",x"87"),
   858 => (x"48",x"72",x"8a",x"0a"),
   859 => (x"4d",x"26",x"87",x"c2"),
   860 => (x"4b",x"26",x"4c",x"26"),
   861 => (x"fd",x"1e",x"4f",x"26"),
   862 => (x"49",x"70",x"87",x"c9"),
   863 => (x"aa",x"f0",x"c0",x"4a"),
   864 => (x"c0",x"87",x"c9",x"04"),
   865 => (x"c3",x"01",x"aa",x"f9"),
   866 => (x"8a",x"f0",x"c0",x"87"),
   867 => (x"04",x"aa",x"c1",x"c1"),
   868 => (x"da",x"c1",x"87",x"c9"),
   869 => (x"87",x"c3",x"01",x"aa"),
   870 => (x"72",x"8a",x"f7",x"c0"),
   871 => (x"0e",x"4f",x"26",x"48"),
   872 => (x"0e",x"5c",x"5b",x"5e"),
   873 => (x"d4",x"ff",x"4a",x"71"),
   874 => (x"c0",x"49",x"72",x"4b"),
   875 => (x"4c",x"70",x"87",x"e7"),
   876 => (x"87",x"c2",x"02",x"9c"),
   877 => (x"d0",x"ff",x"8c",x"c1"),
   878 => (x"c1",x"78",x"c5",x"48"),
   879 => (x"49",x"74",x"7b",x"d5"),
   880 => (x"e9",x"c1",x"31",x"c6"),
   881 => (x"4a",x"bf",x"97",x"da"),
   882 => (x"70",x"b0",x"71",x"48"),
   883 => (x"48",x"d0",x"ff",x"7b"),
   884 => (x"db",x"fe",x"78",x"c4"),
   885 => (x"5b",x"5e",x"0e",x"87"),
   886 => (x"f8",x"0e",x"5d",x"5c"),
   887 => (x"c0",x"4b",x"71",x"86"),
   888 => (x"fc",x"fa",x"c0",x"7e"),
   889 => (x"df",x"49",x"bf",x"97"),
   890 => (x"ee",x"c0",x"05",x"a9"),
   891 => (x"49",x"a3",x"c8",x"87"),
   892 => (x"c1",x"49",x"69",x"97"),
   893 => (x"dd",x"05",x"a9",x"c3"),
   894 => (x"49",x"a3",x"c9",x"87"),
   895 => (x"c1",x"49",x"69",x"97"),
   896 => (x"d1",x"05",x"a9",x"c6"),
   897 => (x"49",x"a3",x"ca",x"87"),
   898 => (x"c1",x"49",x"69",x"97"),
   899 => (x"c5",x"05",x"a9",x"c7"),
   900 => (x"c2",x"48",x"c1",x"87"),
   901 => (x"48",x"c0",x"87",x"e1"),
   902 => (x"fa",x"87",x"dc",x"c2"),
   903 => (x"4c",x"c0",x"87",x"f0"),
   904 => (x"97",x"fc",x"fa",x"c0"),
   905 => (x"a9",x"c0",x"49",x"bf"),
   906 => (x"fb",x"87",x"cf",x"04"),
   907 => (x"84",x"c1",x"87",x"c5"),
   908 => (x"97",x"fc",x"fa",x"c0"),
   909 => (x"06",x"ac",x"49",x"bf"),
   910 => (x"fa",x"c0",x"87",x"f1"),
   911 => (x"02",x"bf",x"97",x"fc"),
   912 => (x"fe",x"f9",x"87",x"cf"),
   913 => (x"99",x"49",x"70",x"87"),
   914 => (x"c0",x"87",x"c6",x"02"),
   915 => (x"f1",x"05",x"a9",x"ec"),
   916 => (x"f9",x"4c",x"c0",x"87"),
   917 => (x"4d",x"70",x"87",x"ed"),
   918 => (x"c8",x"87",x"e8",x"f9"),
   919 => (x"e2",x"f9",x"58",x"a6"),
   920 => (x"c1",x"4a",x"70",x"87"),
   921 => (x"49",x"a3",x"c8",x"84"),
   922 => (x"ad",x"49",x"69",x"97"),
   923 => (x"c0",x"87",x"c7",x"02"),
   924 => (x"c0",x"05",x"ad",x"ff"),
   925 => (x"a3",x"c9",x"87",x"e7"),
   926 => (x"49",x"69",x"97",x"49"),
   927 => (x"02",x"a9",x"66",x"c4"),
   928 => (x"c0",x"48",x"87",x"c7"),
   929 => (x"d4",x"05",x"a8",x"ff"),
   930 => (x"49",x"a3",x"ca",x"87"),
   931 => (x"aa",x"49",x"69",x"97"),
   932 => (x"c0",x"87",x"c6",x"02"),
   933 => (x"c4",x"05",x"aa",x"ff"),
   934 => (x"d0",x"7e",x"c1",x"87"),
   935 => (x"ad",x"ec",x"c0",x"87"),
   936 => (x"c0",x"87",x"c6",x"02"),
   937 => (x"c4",x"05",x"ad",x"fb"),
   938 => (x"c1",x"4c",x"c0",x"87"),
   939 => (x"fe",x"02",x"6e",x"7e"),
   940 => (x"f5",x"f8",x"87",x"e1"),
   941 => (x"f8",x"48",x"74",x"87"),
   942 => (x"87",x"f2",x"fa",x"8e"),
   943 => (x"5b",x"5e",x"0e",x"00"),
   944 => (x"f8",x"0e",x"5d",x"5c"),
   945 => (x"ff",x"4d",x"71",x"86"),
   946 => (x"1e",x"75",x"4b",x"d4"),
   947 => (x"49",x"cc",x"f4",x"c2"),
   948 => (x"c4",x"87",x"ed",x"e4"),
   949 => (x"02",x"98",x"70",x"86"),
   950 => (x"c4",x"87",x"cc",x"c4"),
   951 => (x"e9",x"c1",x"48",x"a6"),
   952 => (x"75",x"78",x"bf",x"dc"),
   953 => (x"87",x"f7",x"fa",x"49"),
   954 => (x"c5",x"48",x"d0",x"ff"),
   955 => (x"7b",x"d6",x"c1",x"78"),
   956 => (x"a2",x"75",x"4a",x"c0"),
   957 => (x"c1",x"7b",x"11",x"49"),
   958 => (x"aa",x"b7",x"cb",x"82"),
   959 => (x"cc",x"87",x"f3",x"04"),
   960 => (x"7b",x"ff",x"c3",x"4a"),
   961 => (x"e0",x"c0",x"82",x"c1"),
   962 => (x"f4",x"04",x"aa",x"b7"),
   963 => (x"48",x"d0",x"ff",x"87"),
   964 => (x"ff",x"c3",x"78",x"c4"),
   965 => (x"c1",x"78",x"c5",x"7b"),
   966 => (x"7b",x"c1",x"7b",x"d3"),
   967 => (x"48",x"66",x"78",x"c4"),
   968 => (x"06",x"a8",x"b7",x"c0"),
   969 => (x"c2",x"87",x"f0",x"c2"),
   970 => (x"4c",x"bf",x"d4",x"f4"),
   971 => (x"74",x"48",x"66",x"c4"),
   972 => (x"58",x"a6",x"c8",x"88"),
   973 => (x"c1",x"02",x"9c",x"74"),
   974 => (x"e7",x"c2",x"87",x"f9"),
   975 => (x"c0",x"c8",x"7e",x"d6"),
   976 => (x"b7",x"c0",x"8c",x"4d"),
   977 => (x"87",x"c6",x"03",x"ac"),
   978 => (x"4d",x"a4",x"c0",x"c8"),
   979 => (x"f4",x"c2",x"4c",x"c0"),
   980 => (x"49",x"bf",x"97",x"c7"),
   981 => (x"d1",x"02",x"99",x"d0"),
   982 => (x"c2",x"1e",x"c0",x"87"),
   983 => (x"e7",x"49",x"cc",x"f4"),
   984 => (x"86",x"c4",x"87",x"d2"),
   985 => (x"c0",x"4a",x"49",x"70"),
   986 => (x"e7",x"c2",x"87",x"ee"),
   987 => (x"f4",x"c2",x"1e",x"d6"),
   988 => (x"ff",x"e6",x"49",x"cc"),
   989 => (x"70",x"86",x"c4",x"87"),
   990 => (x"d0",x"ff",x"4a",x"49"),
   991 => (x"78",x"c5",x"c8",x"48"),
   992 => (x"6e",x"7b",x"d4",x"c1"),
   993 => (x"6e",x"7b",x"bf",x"97"),
   994 => (x"70",x"80",x"c1",x"48"),
   995 => (x"05",x"8d",x"c1",x"7e"),
   996 => (x"ff",x"87",x"f0",x"ff"),
   997 => (x"78",x"c4",x"48",x"d0"),
   998 => (x"c5",x"05",x"9a",x"72"),
   999 => (x"c1",x"48",x"c0",x"87"),
  1000 => (x"1e",x"c1",x"87",x"c7"),
  1001 => (x"49",x"cc",x"f4",x"c2"),
  1002 => (x"c4",x"87",x"ef",x"e4"),
  1003 => (x"05",x"9c",x"74",x"86"),
  1004 => (x"c4",x"87",x"c7",x"fe"),
  1005 => (x"b7",x"c0",x"48",x"66"),
  1006 => (x"87",x"d1",x"06",x"a8"),
  1007 => (x"48",x"cc",x"f4",x"c2"),
  1008 => (x"80",x"d0",x"78",x"c0"),
  1009 => (x"80",x"f4",x"78",x"c0"),
  1010 => (x"bf",x"d8",x"f4",x"c2"),
  1011 => (x"48",x"66",x"c4",x"78"),
  1012 => (x"01",x"a8",x"b7",x"c0"),
  1013 => (x"ff",x"87",x"d0",x"fd"),
  1014 => (x"78",x"c5",x"48",x"d0"),
  1015 => (x"c0",x"7b",x"d3",x"c1"),
  1016 => (x"c1",x"78",x"c4",x"7b"),
  1017 => (x"c0",x"87",x"c2",x"48"),
  1018 => (x"26",x"8e",x"f8",x"48"),
  1019 => (x"26",x"4c",x"26",x"4d"),
  1020 => (x"0e",x"4f",x"26",x"4b"),
  1021 => (x"5d",x"5c",x"5b",x"5e"),
  1022 => (x"4b",x"71",x"1e",x"0e"),
  1023 => (x"ab",x"4d",x"4c",x"c0"),
  1024 => (x"87",x"e8",x"c0",x"04"),
  1025 => (x"1e",x"d5",x"f7",x"c0"),
  1026 => (x"c4",x"02",x"9d",x"75"),
  1027 => (x"c2",x"4a",x"c0",x"87"),
  1028 => (x"72",x"4a",x"c1",x"87"),
  1029 => (x"87",x"f2",x"ea",x"49"),
  1030 => (x"7e",x"70",x"86",x"c4"),
  1031 => (x"05",x"6e",x"84",x"c1"),
  1032 => (x"4c",x"73",x"87",x"c2"),
  1033 => (x"ac",x"73",x"85",x"c1"),
  1034 => (x"87",x"d8",x"ff",x"06"),
  1035 => (x"fe",x"26",x"48",x"6e"),
  1036 => (x"5e",x"0e",x"87",x"f9"),
  1037 => (x"71",x"0e",x"5c",x"5b"),
  1038 => (x"02",x"66",x"cc",x"4b"),
  1039 => (x"4c",x"87",x"e8",x"c0"),
  1040 => (x"02",x"8c",x"f0",x"c0"),
  1041 => (x"74",x"87",x"e8",x"c0"),
  1042 => (x"02",x"8a",x"c1",x"4a"),
  1043 => (x"8a",x"87",x"e0",x"c0"),
  1044 => (x"8a",x"87",x"dc",x"02"),
  1045 => (x"c0",x"87",x"d8",x"02"),
  1046 => (x"c0",x"02",x"8a",x"e0"),
  1047 => (x"8a",x"c1",x"87",x"e5"),
  1048 => (x"87",x"e7",x"c0",x"02"),
  1049 => (x"73",x"87",x"ea",x"c0"),
  1050 => (x"87",x"d1",x"f9",x"49"),
  1051 => (x"74",x"87",x"e2",x"c0"),
  1052 => (x"c1",x"49",x"c0",x"1e"),
  1053 => (x"74",x"87",x"d2",x"e0"),
  1054 => (x"c1",x"49",x"73",x"1e"),
  1055 => (x"c8",x"87",x"ca",x"e0"),
  1056 => (x"73",x"87",x"ce",x"86"),
  1057 => (x"f5",x"e2",x"c1",x"49"),
  1058 => (x"73",x"87",x"c6",x"87"),
  1059 => (x"e5",x"e3",x"c1",x"49"),
  1060 => (x"87",x"d9",x"fd",x"87"),
  1061 => (x"5c",x"5b",x"5e",x"0e"),
  1062 => (x"71",x"1e",x"0e",x"5d"),
  1063 => (x"91",x"de",x"49",x"4c"),
  1064 => (x"4d",x"f4",x"f4",x"c2"),
  1065 => (x"6d",x"97",x"85",x"71"),
  1066 => (x"87",x"de",x"c1",x"02"),
  1067 => (x"bf",x"e0",x"f4",x"c2"),
  1068 => (x"72",x"82",x"74",x"4a"),
  1069 => (x"87",x"fb",x"fc",x"49"),
  1070 => (x"98",x"48",x"7e",x"70"),
  1071 => (x"87",x"f2",x"c0",x"02"),
  1072 => (x"4b",x"e8",x"f4",x"c2"),
  1073 => (x"49",x"cb",x"4a",x"70"),
  1074 => (x"87",x"db",x"ff",x"fe"),
  1075 => (x"93",x"cb",x"4b",x"74"),
  1076 => (x"83",x"d1",x"ea",x"c1"),
  1077 => (x"c4",x"c1",x"83",x"c4"),
  1078 => (x"49",x"74",x"7b",x"ce"),
  1079 => (x"87",x"d2",x"c6",x"c1"),
  1080 => (x"e9",x"c1",x"7b",x"75"),
  1081 => (x"49",x"bf",x"97",x"db"),
  1082 => (x"e8",x"f4",x"c2",x"1e"),
  1083 => (x"87",x"c2",x"fd",x"49"),
  1084 => (x"49",x"74",x"86",x"c4"),
  1085 => (x"87",x"fa",x"c5",x"c1"),
  1086 => (x"c7",x"c1",x"49",x"c0"),
  1087 => (x"f4",x"c2",x"87",x"d9"),
  1088 => (x"78",x"c0",x"48",x"c8"),
  1089 => (x"e0",x"c0",x"49",x"c1"),
  1090 => (x"fb",x"26",x"87",x"ff"),
  1091 => (x"6f",x"4c",x"87",x"dd"),
  1092 => (x"6e",x"69",x"64",x"61"),
  1093 => (x"2e",x"2e",x"2e",x"67"),
  1094 => (x"5b",x"5e",x"0e",x"00"),
  1095 => (x"4b",x"71",x"0e",x"5c"),
  1096 => (x"e0",x"f4",x"c2",x"4a"),
  1097 => (x"49",x"72",x"82",x"bf"),
  1098 => (x"70",x"87",x"c8",x"fb"),
  1099 => (x"c4",x"02",x"9c",x"4c"),
  1100 => (x"dd",x"e5",x"49",x"87"),
  1101 => (x"e0",x"f4",x"c2",x"87"),
  1102 => (x"c1",x"78",x"c0",x"48"),
  1103 => (x"c8",x"e0",x"c0",x"49"),
  1104 => (x"87",x"e9",x"fa",x"87"),
  1105 => (x"5c",x"5b",x"5e",x"0e"),
  1106 => (x"86",x"f4",x"0e",x"5d"),
  1107 => (x"4d",x"d6",x"e7",x"c2"),
  1108 => (x"a6",x"c4",x"4c",x"c0"),
  1109 => (x"c2",x"78",x"c0",x"48"),
  1110 => (x"49",x"bf",x"e0",x"f4"),
  1111 => (x"c1",x"06",x"a9",x"c0"),
  1112 => (x"e7",x"c2",x"87",x"c1"),
  1113 => (x"02",x"98",x"48",x"d6"),
  1114 => (x"c0",x"87",x"f8",x"c0"),
  1115 => (x"c8",x"1e",x"d5",x"f7"),
  1116 => (x"87",x"c7",x"02",x"66"),
  1117 => (x"c0",x"48",x"a6",x"c4"),
  1118 => (x"c4",x"87",x"c5",x"78"),
  1119 => (x"78",x"c1",x"48",x"a6"),
  1120 => (x"e5",x"49",x"66",x"c4"),
  1121 => (x"86",x"c4",x"87",x"c4"),
  1122 => (x"84",x"c1",x"4d",x"70"),
  1123 => (x"c1",x"48",x"66",x"c4"),
  1124 => (x"58",x"a6",x"c8",x"80"),
  1125 => (x"bf",x"e0",x"f4",x"c2"),
  1126 => (x"c6",x"03",x"ac",x"49"),
  1127 => (x"05",x"9d",x"75",x"87"),
  1128 => (x"c0",x"87",x"c8",x"ff"),
  1129 => (x"02",x"9d",x"75",x"4c"),
  1130 => (x"c0",x"87",x"e0",x"c3"),
  1131 => (x"c8",x"1e",x"d5",x"f7"),
  1132 => (x"87",x"c7",x"02",x"66"),
  1133 => (x"c0",x"48",x"a6",x"cc"),
  1134 => (x"cc",x"87",x"c5",x"78"),
  1135 => (x"78",x"c1",x"48",x"a6"),
  1136 => (x"e4",x"49",x"66",x"cc"),
  1137 => (x"86",x"c4",x"87",x"c4"),
  1138 => (x"98",x"48",x"7e",x"70"),
  1139 => (x"87",x"e8",x"c2",x"02"),
  1140 => (x"97",x"81",x"cb",x"49"),
  1141 => (x"99",x"d0",x"49",x"69"),
  1142 => (x"87",x"d6",x"c1",x"02"),
  1143 => (x"4a",x"d9",x"c4",x"c1"),
  1144 => (x"91",x"cb",x"49",x"74"),
  1145 => (x"81",x"d1",x"ea",x"c1"),
  1146 => (x"81",x"c8",x"79",x"72"),
  1147 => (x"74",x"51",x"ff",x"c3"),
  1148 => (x"c2",x"91",x"de",x"49"),
  1149 => (x"71",x"4d",x"f4",x"f4"),
  1150 => (x"97",x"c1",x"c2",x"85"),
  1151 => (x"49",x"a5",x"c1",x"7d"),
  1152 => (x"c2",x"51",x"e0",x"c0"),
  1153 => (x"bf",x"97",x"e6",x"ef"),
  1154 => (x"c1",x"87",x"d2",x"02"),
  1155 => (x"4b",x"a5",x"c2",x"84"),
  1156 => (x"4a",x"e6",x"ef",x"c2"),
  1157 => (x"fa",x"fe",x"49",x"db"),
  1158 => (x"db",x"c1",x"87",x"cd"),
  1159 => (x"49",x"a5",x"cd",x"87"),
  1160 => (x"84",x"c1",x"51",x"c0"),
  1161 => (x"6e",x"4b",x"a5",x"c2"),
  1162 => (x"fe",x"49",x"cb",x"4a"),
  1163 => (x"c1",x"87",x"f8",x"f9"),
  1164 => (x"c2",x"c1",x"87",x"c6"),
  1165 => (x"49",x"74",x"4a",x"d4"),
  1166 => (x"ea",x"c1",x"91",x"cb"),
  1167 => (x"79",x"72",x"81",x"d1"),
  1168 => (x"97",x"e6",x"ef",x"c2"),
  1169 => (x"87",x"d8",x"02",x"bf"),
  1170 => (x"91",x"de",x"49",x"74"),
  1171 => (x"f4",x"c2",x"84",x"c1"),
  1172 => (x"83",x"71",x"4b",x"f4"),
  1173 => (x"4a",x"e6",x"ef",x"c2"),
  1174 => (x"f9",x"fe",x"49",x"dd"),
  1175 => (x"87",x"d8",x"87",x"c9"),
  1176 => (x"93",x"de",x"4b",x"74"),
  1177 => (x"83",x"f4",x"f4",x"c2"),
  1178 => (x"c0",x"49",x"a3",x"cb"),
  1179 => (x"73",x"84",x"c1",x"51"),
  1180 => (x"49",x"cb",x"4a",x"6e"),
  1181 => (x"87",x"ef",x"f8",x"fe"),
  1182 => (x"c1",x"48",x"66",x"c4"),
  1183 => (x"58",x"a6",x"c8",x"80"),
  1184 => (x"c0",x"03",x"ac",x"c7"),
  1185 => (x"05",x"6e",x"87",x"c5"),
  1186 => (x"74",x"87",x"e0",x"fc"),
  1187 => (x"f5",x"8e",x"f4",x"48"),
  1188 => (x"73",x"1e",x"87",x"d9"),
  1189 => (x"49",x"4b",x"71",x"1e"),
  1190 => (x"ea",x"c1",x"91",x"cb"),
  1191 => (x"a1",x"c8",x"81",x"d1"),
  1192 => (x"da",x"e9",x"c1",x"4a"),
  1193 => (x"c9",x"50",x"12",x"48"),
  1194 => (x"fa",x"c0",x"4a",x"a1"),
  1195 => (x"50",x"12",x"48",x"fc"),
  1196 => (x"e9",x"c1",x"81",x"ca"),
  1197 => (x"50",x"11",x"48",x"db"),
  1198 => (x"97",x"db",x"e9",x"c1"),
  1199 => (x"c0",x"1e",x"49",x"bf"),
  1200 => (x"87",x"ee",x"f5",x"49"),
  1201 => (x"48",x"c8",x"f4",x"c2"),
  1202 => (x"49",x"c1",x"78",x"de"),
  1203 => (x"26",x"87",x"fa",x"d9"),
  1204 => (x"1e",x"87",x"dc",x"f4"),
  1205 => (x"cb",x"49",x"4a",x"71"),
  1206 => (x"d1",x"ea",x"c1",x"91"),
  1207 => (x"11",x"81",x"c8",x"81"),
  1208 => (x"cc",x"f4",x"c2",x"48"),
  1209 => (x"e0",x"f4",x"c2",x"58"),
  1210 => (x"c1",x"78",x"c0",x"48"),
  1211 => (x"87",x"d9",x"d9",x"49"),
  1212 => (x"c0",x"1e",x"4f",x"26"),
  1213 => (x"de",x"ff",x"c0",x"49"),
  1214 => (x"1e",x"4f",x"26",x"87"),
  1215 => (x"d2",x"02",x"99",x"71"),
  1216 => (x"e6",x"eb",x"c1",x"87"),
  1217 => (x"f7",x"50",x"c0",x"48"),
  1218 => (x"d3",x"cb",x"c1",x"80"),
  1219 => (x"ff",x"e9",x"c1",x"40"),
  1220 => (x"c1",x"87",x"ce",x"78"),
  1221 => (x"c1",x"48",x"e2",x"eb"),
  1222 => (x"fc",x"78",x"e0",x"e9"),
  1223 => (x"f2",x"cb",x"c1",x"80"),
  1224 => (x"0e",x"4f",x"26",x"78"),
  1225 => (x"5d",x"5c",x"5b",x"5e"),
  1226 => (x"71",x"86",x"f4",x"0e"),
  1227 => (x"91",x"cb",x"49",x"4d"),
  1228 => (x"81",x"d1",x"ea",x"c1"),
  1229 => (x"ca",x"4a",x"a1",x"c8"),
  1230 => (x"a6",x"c4",x"7e",x"a1"),
  1231 => (x"d0",x"f8",x"c2",x"48"),
  1232 => (x"97",x"6e",x"78",x"bf"),
  1233 => (x"66",x"c4",x"4b",x"bf"),
  1234 => (x"70",x"28",x"73",x"48"),
  1235 => (x"48",x"12",x"4c",x"4b"),
  1236 => (x"70",x"58",x"a6",x"cc"),
  1237 => (x"c9",x"84",x"c1",x"9c"),
  1238 => (x"49",x"69",x"97",x"81"),
  1239 => (x"c2",x"04",x"ac",x"b7"),
  1240 => (x"6e",x"4c",x"c0",x"87"),
  1241 => (x"c8",x"4a",x"bf",x"97"),
  1242 => (x"31",x"72",x"49",x"66"),
  1243 => (x"66",x"c4",x"b9",x"ff"),
  1244 => (x"72",x"48",x"74",x"99"),
  1245 => (x"48",x"4a",x"70",x"30"),
  1246 => (x"f8",x"c2",x"b0",x"71"),
  1247 => (x"e9",x"c0",x"58",x"d4"),
  1248 => (x"49",x"c0",x"87",x"f0"),
  1249 => (x"75",x"87",x"c2",x"d7"),
  1250 => (x"e5",x"fb",x"c0",x"49"),
  1251 => (x"f1",x"8e",x"f4",x"87"),
  1252 => (x"73",x"1e",x"87",x"d9"),
  1253 => (x"49",x"4b",x"71",x"1e"),
  1254 => (x"73",x"87",x"c8",x"fe"),
  1255 => (x"87",x"c3",x"fe",x"49"),
  1256 => (x"1e",x"87",x"cc",x"f1"),
  1257 => (x"4b",x"71",x"1e",x"73"),
  1258 => (x"02",x"4a",x"a3",x"c6"),
  1259 => (x"8a",x"c1",x"87",x"dc"),
  1260 => (x"87",x"e4",x"c0",x"02"),
  1261 => (x"e8",x"c1",x"02",x"8a"),
  1262 => (x"c1",x"02",x"8a",x"87"),
  1263 => (x"02",x"8a",x"87",x"ca"),
  1264 => (x"8a",x"87",x"ef",x"c0"),
  1265 => (x"c1",x"87",x"d9",x"02"),
  1266 => (x"f4",x"c2",x"87",x"e9"),
  1267 => (x"78",x"df",x"48",x"c8"),
  1268 => (x"f4",x"d5",x"49",x"c1"),
  1269 => (x"87",x"e6",x"c1",x"87"),
  1270 => (x"f6",x"fb",x"49",x"c7"),
  1271 => (x"87",x"de",x"c1",x"87"),
  1272 => (x"bf",x"e0",x"f4",x"c2"),
  1273 => (x"87",x"cb",x"c1",x"02"),
  1274 => (x"c2",x"88",x"c1",x"48"),
  1275 => (x"c1",x"58",x"e4",x"f4"),
  1276 => (x"f4",x"c2",x"87",x"c1"),
  1277 => (x"c0",x"02",x"bf",x"e4"),
  1278 => (x"f4",x"c2",x"87",x"f9"),
  1279 => (x"c1",x"48",x"bf",x"e0"),
  1280 => (x"e4",x"f4",x"c2",x"80"),
  1281 => (x"87",x"eb",x"c0",x"58"),
  1282 => (x"bf",x"e0",x"f4",x"c2"),
  1283 => (x"c2",x"89",x"c6",x"49"),
  1284 => (x"c0",x"59",x"e4",x"f4"),
  1285 => (x"da",x"03",x"a9",x"b7"),
  1286 => (x"e0",x"f4",x"c2",x"87"),
  1287 => (x"d2",x"78",x"c0",x"48"),
  1288 => (x"e4",x"f4",x"c2",x"87"),
  1289 => (x"87",x"cb",x"02",x"bf"),
  1290 => (x"bf",x"e0",x"f4",x"c2"),
  1291 => (x"c2",x"80",x"c6",x"48"),
  1292 => (x"c0",x"58",x"e4",x"f4"),
  1293 => (x"87",x"d1",x"d4",x"49"),
  1294 => (x"f8",x"c0",x"49",x"73"),
  1295 => (x"ee",x"ee",x"87",x"f4"),
  1296 => (x"5b",x"5e",x"0e",x"87"),
  1297 => (x"ff",x"0e",x"5d",x"5c"),
  1298 => (x"a6",x"dc",x"86",x"d0"),
  1299 => (x"cc",x"4d",x"c0",x"59"),
  1300 => (x"c4",x"c1",x"48",x"a6"),
  1301 => (x"80",x"c4",x"78",x"66"),
  1302 => (x"80",x"c4",x"78",x"c1"),
  1303 => (x"f4",x"c2",x"78",x"c1"),
  1304 => (x"78",x"c1",x"48",x"e4"),
  1305 => (x"bf",x"c8",x"f4",x"c2"),
  1306 => (x"de",x"48",x"6e",x"7e"),
  1307 => (x"87",x"c9",x"05",x"a8"),
  1308 => (x"70",x"87",x"d1",x"f3"),
  1309 => (x"f9",x"d1",x"4d",x"49"),
  1310 => (x"df",x"48",x"6e",x"87"),
  1311 => (x"eb",x"c1",x"05",x"a8"),
  1312 => (x"66",x"c0",x"c1",x"87"),
  1313 => (x"69",x"81",x"c4",x"49"),
  1314 => (x"dd",x"e4",x"c1",x"7e"),
  1315 => (x"d0",x"49",x"6e",x"48"),
  1316 => (x"41",x"20",x"4a",x"a1"),
  1317 => (x"f9",x"05",x"aa",x"71"),
  1318 => (x"d2",x"ca",x"c1",x"87"),
  1319 => (x"66",x"c0",x"c1",x"4a"),
  1320 => (x"c1",x"0a",x"7a",x"0a"),
  1321 => (x"c9",x"49",x"66",x"c0"),
  1322 => (x"c1",x"51",x"df",x"81"),
  1323 => (x"ca",x"49",x"66",x"c0"),
  1324 => (x"51",x"d3",x"c1",x"81"),
  1325 => (x"49",x"66",x"c0",x"c1"),
  1326 => (x"a1",x"c4",x"81",x"cb"),
  1327 => (x"48",x"a6",x"c4",x"4b"),
  1328 => (x"1e",x"71",x"78",x"6b"),
  1329 => (x"e4",x"c1",x"1e",x"72"),
  1330 => (x"66",x"cc",x"48",x"ed"),
  1331 => (x"4a",x"a1",x"d0",x"49"),
  1332 => (x"aa",x"71",x"41",x"20"),
  1333 => (x"26",x"87",x"f9",x"05"),
  1334 => (x"72",x"49",x"26",x"4a"),
  1335 => (x"4a",x"a1",x"c9",x"79"),
  1336 => (x"81",x"ca",x"52",x"df"),
  1337 => (x"c2",x"51",x"d4",x"c1"),
  1338 => (x"87",x"c6",x"d0",x"4d"),
  1339 => (x"87",x"de",x"df",x"ff"),
  1340 => (x"ff",x"87",x"c0",x"e0"),
  1341 => (x"70",x"87",x"cc",x"df"),
  1342 => (x"ac",x"fb",x"c0",x"4c"),
  1343 => (x"87",x"fa",x"c1",x"02"),
  1344 => (x"c1",x"05",x"66",x"d8"),
  1345 => (x"c0",x"c1",x"87",x"eb"),
  1346 => (x"82",x"c4",x"4a",x"66"),
  1347 => (x"1e",x"72",x"7e",x"6a"),
  1348 => (x"48",x"fd",x"e4",x"c1"),
  1349 => (x"c8",x"49",x"66",x"c4"),
  1350 => (x"41",x"20",x"4a",x"a1"),
  1351 => (x"f9",x"05",x"aa",x"71"),
  1352 => (x"26",x"51",x"10",x"87"),
  1353 => (x"66",x"c0",x"c1",x"4a"),
  1354 => (x"d2",x"ca",x"c1",x"48"),
  1355 => (x"c7",x"49",x"6a",x"78"),
  1356 => (x"c1",x"51",x"74",x"81"),
  1357 => (x"c8",x"49",x"66",x"c0"),
  1358 => (x"c1",x"51",x"c1",x"81"),
  1359 => (x"c9",x"49",x"66",x"c0"),
  1360 => (x"c1",x"51",x"c0",x"81"),
  1361 => (x"ca",x"49",x"66",x"c0"),
  1362 => (x"c1",x"51",x"c0",x"81"),
  1363 => (x"6a",x"1e",x"d8",x"1e"),
  1364 => (x"ff",x"81",x"c8",x"49"),
  1365 => (x"c8",x"87",x"f0",x"de"),
  1366 => (x"66",x"c4",x"c1",x"86"),
  1367 => (x"01",x"a8",x"c0",x"48"),
  1368 => (x"4d",x"c1",x"87",x"c4"),
  1369 => (x"c4",x"c1",x"87",x"cf"),
  1370 => (x"88",x"c1",x"48",x"66"),
  1371 => (x"c4",x"58",x"a6",x"d0"),
  1372 => (x"fe",x"dd",x"ff",x"87"),
  1373 => (x"48",x"a6",x"d0",x"87"),
  1374 => (x"a6",x"cc",x"78",x"c2"),
  1375 => (x"02",x"9c",x"74",x"5d"),
  1376 => (x"cc",x"87",x"e8",x"cd"),
  1377 => (x"c8",x"c1",x"5d",x"a6"),
  1378 => (x"cd",x"03",x"ad",x"66"),
  1379 => (x"a6",x"dc",x"87",x"dd"),
  1380 => (x"e8",x"78",x"c0",x"48"),
  1381 => (x"ff",x"78",x"c0",x"80"),
  1382 => (x"70",x"87",x"e8",x"dc"),
  1383 => (x"ac",x"d0",x"c1",x"4c"),
  1384 => (x"87",x"db",x"c2",x"05"),
  1385 => (x"ff",x"7e",x"66",x"c4"),
  1386 => (x"70",x"87",x"cb",x"df"),
  1387 => (x"59",x"a6",x"c8",x"49"),
  1388 => (x"87",x"cf",x"dc",x"ff"),
  1389 => (x"ec",x"c0",x"4c",x"70"),
  1390 => (x"ed",x"c1",x"05",x"ac"),
  1391 => (x"49",x"66",x"c8",x"87"),
  1392 => (x"c0",x"c1",x"91",x"cb"),
  1393 => (x"a1",x"c4",x"81",x"66"),
  1394 => (x"c8",x"4d",x"6a",x"4a"),
  1395 => (x"66",x"c4",x"4a",x"a1"),
  1396 => (x"d3",x"cb",x"c1",x"52"),
  1397 => (x"ea",x"db",x"ff",x"79"),
  1398 => (x"9c",x"4c",x"70",x"87"),
  1399 => (x"c0",x"87",x"d9",x"02"),
  1400 => (x"d3",x"02",x"ac",x"fb"),
  1401 => (x"ff",x"55",x"74",x"87"),
  1402 => (x"70",x"87",x"d8",x"db"),
  1403 => (x"c7",x"02",x"9c",x"4c"),
  1404 => (x"ac",x"fb",x"c0",x"87"),
  1405 => (x"87",x"ed",x"ff",x"05"),
  1406 => (x"c2",x"55",x"e0",x"c0"),
  1407 => (x"97",x"c0",x"55",x"c1"),
  1408 => (x"49",x"66",x"d8",x"7d"),
  1409 => (x"db",x"05",x"a9",x"6e"),
  1410 => (x"48",x"66",x"c8",x"87"),
  1411 => (x"04",x"a8",x"66",x"cc"),
  1412 => (x"66",x"c8",x"87",x"ca"),
  1413 => (x"cc",x"80",x"c1",x"48"),
  1414 => (x"87",x"c8",x"58",x"a6"),
  1415 => (x"c1",x"48",x"66",x"cc"),
  1416 => (x"58",x"a6",x"d0",x"88"),
  1417 => (x"87",x"db",x"da",x"ff"),
  1418 => (x"d0",x"c1",x"4c",x"70"),
  1419 => (x"87",x"c8",x"05",x"ac"),
  1420 => (x"c1",x"48",x"66",x"d4"),
  1421 => (x"58",x"a6",x"d8",x"80"),
  1422 => (x"02",x"ac",x"d0",x"c1"),
  1423 => (x"c0",x"87",x"e5",x"fd"),
  1424 => (x"d8",x"48",x"a6",x"e0"),
  1425 => (x"66",x"c4",x"78",x"66"),
  1426 => (x"66",x"e0",x"c0",x"48"),
  1427 => (x"ec",x"c9",x"05",x"a8"),
  1428 => (x"a6",x"e4",x"c0",x"87"),
  1429 => (x"74",x"78",x"c0",x"48"),
  1430 => (x"88",x"fb",x"c0",x"48"),
  1431 => (x"98",x"48",x"7e",x"70"),
  1432 => (x"87",x"ee",x"c9",x"02"),
  1433 => (x"70",x"88",x"cb",x"48"),
  1434 => (x"02",x"98",x"48",x"7e"),
  1435 => (x"48",x"87",x"ce",x"c1"),
  1436 => (x"7e",x"70",x"88",x"c9"),
  1437 => (x"c4",x"02",x"98",x"48"),
  1438 => (x"c4",x"48",x"87",x"c2"),
  1439 => (x"48",x"7e",x"70",x"88"),
  1440 => (x"87",x"ce",x"02",x"98"),
  1441 => (x"70",x"88",x"c1",x"48"),
  1442 => (x"02",x"98",x"48",x"7e"),
  1443 => (x"c8",x"87",x"ed",x"c3"),
  1444 => (x"a6",x"dc",x"87",x"e2"),
  1445 => (x"78",x"f0",x"c0",x"48"),
  1446 => (x"87",x"e7",x"d8",x"ff"),
  1447 => (x"ec",x"c0",x"4c",x"70"),
  1448 => (x"c4",x"c0",x"02",x"ac"),
  1449 => (x"a6",x"e0",x"c0",x"87"),
  1450 => (x"ac",x"ec",x"c0",x"5c"),
  1451 => (x"87",x"cd",x"c0",x"02"),
  1452 => (x"87",x"cf",x"d8",x"ff"),
  1453 => (x"ec",x"c0",x"4c",x"70"),
  1454 => (x"f3",x"ff",x"05",x"ac"),
  1455 => (x"ac",x"ec",x"c0",x"87"),
  1456 => (x"87",x"c4",x"c0",x"02"),
  1457 => (x"87",x"fb",x"d7",x"ff"),
  1458 => (x"1e",x"ca",x"1e",x"c0"),
  1459 => (x"cb",x"49",x"66",x"d0"),
  1460 => (x"66",x"c8",x"c1",x"91"),
  1461 => (x"cc",x"80",x"71",x"48"),
  1462 => (x"66",x"c8",x"58",x"a6"),
  1463 => (x"d0",x"80",x"c4",x"48"),
  1464 => (x"66",x"cc",x"58",x"a6"),
  1465 => (x"d8",x"ff",x"49",x"bf"),
  1466 => (x"1e",x"c1",x"87",x"dd"),
  1467 => (x"66",x"d4",x"1e",x"de"),
  1468 => (x"d8",x"ff",x"49",x"bf"),
  1469 => (x"86",x"d0",x"87",x"d1"),
  1470 => (x"09",x"c0",x"49",x"70"),
  1471 => (x"a6",x"ec",x"c0",x"89"),
  1472 => (x"66",x"e8",x"c0",x"59"),
  1473 => (x"06",x"a8",x"c0",x"48"),
  1474 => (x"c0",x"87",x"ee",x"c0"),
  1475 => (x"dd",x"48",x"66",x"e8"),
  1476 => (x"e4",x"c0",x"03",x"a8"),
  1477 => (x"bf",x"66",x"c4",x"87"),
  1478 => (x"66",x"e8",x"c0",x"49"),
  1479 => (x"51",x"e0",x"c0",x"81"),
  1480 => (x"49",x"66",x"e8",x"c0"),
  1481 => (x"66",x"c4",x"81",x"c1"),
  1482 => (x"c1",x"c2",x"81",x"bf"),
  1483 => (x"66",x"e8",x"c0",x"51"),
  1484 => (x"c4",x"81",x"c2",x"49"),
  1485 => (x"c0",x"81",x"bf",x"66"),
  1486 => (x"c1",x"48",x"6e",x"51"),
  1487 => (x"6e",x"78",x"d2",x"ca"),
  1488 => (x"d0",x"81",x"c8",x"49"),
  1489 => (x"49",x"6e",x"51",x"66"),
  1490 => (x"66",x"d4",x"81",x"c9"),
  1491 => (x"ca",x"49",x"6e",x"51"),
  1492 => (x"51",x"66",x"dc",x"81"),
  1493 => (x"c1",x"48",x"66",x"d0"),
  1494 => (x"58",x"a6",x"d4",x"80"),
  1495 => (x"cc",x"48",x"66",x"c8"),
  1496 => (x"c0",x"04",x"a8",x"66"),
  1497 => (x"66",x"c8",x"87",x"cb"),
  1498 => (x"cc",x"80",x"c1",x"48"),
  1499 => (x"e1",x"c5",x"58",x"a6"),
  1500 => (x"48",x"66",x"cc",x"87"),
  1501 => (x"a6",x"d0",x"88",x"c1"),
  1502 => (x"87",x"d6",x"c5",x"58"),
  1503 => (x"87",x"f6",x"d7",x"ff"),
  1504 => (x"ec",x"c0",x"49",x"70"),
  1505 => (x"d7",x"ff",x"59",x"a6"),
  1506 => (x"49",x"70",x"87",x"ec"),
  1507 => (x"59",x"a6",x"e0",x"c0"),
  1508 => (x"c0",x"48",x"66",x"dc"),
  1509 => (x"c0",x"05",x"a8",x"ec"),
  1510 => (x"a6",x"dc",x"87",x"ca"),
  1511 => (x"66",x"e8",x"c0",x"48"),
  1512 => (x"87",x"c4",x"c0",x"78"),
  1513 => (x"87",x"db",x"d4",x"ff"),
  1514 => (x"cb",x"49",x"66",x"c8"),
  1515 => (x"66",x"c0",x"c1",x"91"),
  1516 => (x"70",x"80",x"71",x"48"),
  1517 => (x"82",x"c8",x"4a",x"7e"),
  1518 => (x"81",x"ca",x"49",x"6e"),
  1519 => (x"51",x"66",x"e8",x"c0"),
  1520 => (x"c1",x"49",x"66",x"dc"),
  1521 => (x"66",x"e8",x"c0",x"81"),
  1522 => (x"71",x"48",x"c1",x"89"),
  1523 => (x"c1",x"49",x"70",x"30"),
  1524 => (x"7a",x"97",x"71",x"89"),
  1525 => (x"bf",x"d0",x"f8",x"c2"),
  1526 => (x"66",x"e8",x"c0",x"49"),
  1527 => (x"4a",x"6a",x"97",x"29"),
  1528 => (x"c0",x"98",x"71",x"48"),
  1529 => (x"6e",x"58",x"a6",x"f0"),
  1530 => (x"69",x"81",x"c4",x"49"),
  1531 => (x"66",x"e0",x"c0",x"4d"),
  1532 => (x"a8",x"66",x"c4",x"48"),
  1533 => (x"87",x"c8",x"c0",x"02"),
  1534 => (x"c0",x"48",x"a6",x"c4"),
  1535 => (x"87",x"c5",x"c0",x"78"),
  1536 => (x"c1",x"48",x"a6",x"c4"),
  1537 => (x"1e",x"66",x"c4",x"78"),
  1538 => (x"75",x"1e",x"e0",x"c0"),
  1539 => (x"f6",x"d3",x"ff",x"49"),
  1540 => (x"70",x"86",x"c8",x"87"),
  1541 => (x"ac",x"b7",x"c0",x"4c"),
  1542 => (x"87",x"d4",x"c1",x"06"),
  1543 => (x"e0",x"c0",x"85",x"74"),
  1544 => (x"75",x"89",x"74",x"49"),
  1545 => (x"c6",x"e5",x"c1",x"4b"),
  1546 => (x"e1",x"fe",x"71",x"4a"),
  1547 => (x"85",x"c2",x"87",x"f9"),
  1548 => (x"48",x"66",x"e4",x"c0"),
  1549 => (x"e8",x"c0",x"80",x"c1"),
  1550 => (x"ec",x"c0",x"58",x"a6"),
  1551 => (x"81",x"c1",x"49",x"66"),
  1552 => (x"c0",x"02",x"a9",x"70"),
  1553 => (x"a6",x"c4",x"87",x"c8"),
  1554 => (x"c0",x"78",x"c0",x"48"),
  1555 => (x"a6",x"c4",x"87",x"c5"),
  1556 => (x"c4",x"78",x"c1",x"48"),
  1557 => (x"a4",x"c2",x"1e",x"66"),
  1558 => (x"48",x"e0",x"c0",x"49"),
  1559 => (x"49",x"70",x"88",x"71"),
  1560 => (x"ff",x"49",x"75",x"1e"),
  1561 => (x"c8",x"87",x"e0",x"d2"),
  1562 => (x"a8",x"b7",x"c0",x"86"),
  1563 => (x"87",x"c0",x"ff",x"01"),
  1564 => (x"02",x"66",x"e4",x"c0"),
  1565 => (x"6e",x"87",x"d1",x"c0"),
  1566 => (x"c0",x"81",x"c9",x"49"),
  1567 => (x"6e",x"51",x"66",x"e4"),
  1568 => (x"e3",x"cc",x"c1",x"48"),
  1569 => (x"87",x"cc",x"c0",x"78"),
  1570 => (x"81",x"c9",x"49",x"6e"),
  1571 => (x"48",x"6e",x"51",x"c2"),
  1572 => (x"78",x"d2",x"ce",x"c1"),
  1573 => (x"cc",x"48",x"66",x"c8"),
  1574 => (x"c0",x"04",x"a8",x"66"),
  1575 => (x"66",x"c8",x"87",x"cb"),
  1576 => (x"cc",x"80",x"c1",x"48"),
  1577 => (x"e9",x"c0",x"58",x"a6"),
  1578 => (x"48",x"66",x"cc",x"87"),
  1579 => (x"a6",x"d0",x"88",x"c1"),
  1580 => (x"87",x"de",x"c0",x"58"),
  1581 => (x"87",x"fb",x"d0",x"ff"),
  1582 => (x"d5",x"c0",x"4c",x"70"),
  1583 => (x"ac",x"c6",x"c1",x"87"),
  1584 => (x"87",x"c8",x"c0",x"05"),
  1585 => (x"c1",x"48",x"66",x"d0"),
  1586 => (x"58",x"a6",x"d4",x"80"),
  1587 => (x"87",x"e3",x"d0",x"ff"),
  1588 => (x"66",x"d4",x"4c",x"70"),
  1589 => (x"d8",x"80",x"c1",x"48"),
  1590 => (x"9c",x"74",x"58",x"a6"),
  1591 => (x"87",x"cb",x"c0",x"02"),
  1592 => (x"c1",x"48",x"66",x"c8"),
  1593 => (x"04",x"a8",x"66",x"c8"),
  1594 => (x"c8",x"87",x"e3",x"f2"),
  1595 => (x"cf",x"ff",x"4d",x"66"),
  1596 => (x"ad",x"c7",x"87",x"f8"),
  1597 => (x"87",x"de",x"c0",x"03"),
  1598 => (x"48",x"e4",x"f4",x"c2"),
  1599 => (x"49",x"75",x"78",x"c0"),
  1600 => (x"c0",x"c1",x"91",x"cb"),
  1601 => (x"a1",x"c4",x"81",x"66"),
  1602 => (x"c0",x"4a",x"6a",x"4a"),
  1603 => (x"85",x"c1",x"79",x"52"),
  1604 => (x"ff",x"04",x"ad",x"c7"),
  1605 => (x"d0",x"ff",x"87",x"e2"),
  1606 => (x"ce",x"db",x"ff",x"8e"),
  1607 => (x"61",x"6f",x"4c",x"87"),
  1608 => (x"65",x"53",x"20",x"64"),
  1609 => (x"6e",x"69",x"74",x"74"),
  1610 => (x"81",x"20",x"73",x"67"),
  1611 => (x"76",x"61",x"53",x"00"),
  1612 => (x"65",x"53",x"20",x"65"),
  1613 => (x"6e",x"69",x"74",x"74"),
  1614 => (x"81",x"20",x"73",x"67"),
  1615 => (x"61",x"6f",x"4c",x"00"),
  1616 => (x"2e",x"2a",x"20",x"64"),
  1617 => (x"20",x"3a",x"00",x"20"),
  1618 => (x"1e",x"73",x"1e",x"00"),
  1619 => (x"02",x"9b",x"4b",x"71"),
  1620 => (x"f4",x"c2",x"87",x"c6"),
  1621 => (x"78",x"c0",x"48",x"e0"),
  1622 => (x"f4",x"c2",x"1e",x"c7"),
  1623 => (x"1e",x"49",x"bf",x"e0"),
  1624 => (x"1e",x"d1",x"ea",x"c1"),
  1625 => (x"bf",x"c8",x"f4",x"c2"),
  1626 => (x"87",x"d5",x"eb",x"49"),
  1627 => (x"f4",x"c2",x"86",x"cc"),
  1628 => (x"e6",x"49",x"bf",x"c8"),
  1629 => (x"9b",x"73",x"87",x"c5"),
  1630 => (x"c1",x"87",x"c8",x"02"),
  1631 => (x"c0",x"49",x"d1",x"ea"),
  1632 => (x"ff",x"87",x"c1",x"e5"),
  1633 => (x"1e",x"87",x"e8",x"d9"),
  1634 => (x"4b",x"c0",x"1e",x"73"),
  1635 => (x"49",x"f2",x"e6",x"c1"),
  1636 => (x"87",x"ea",x"fe",x"c0"),
  1637 => (x"48",x"da",x"e9",x"c1"),
  1638 => (x"eb",x"c1",x"50",x"c0"),
  1639 => (x"ff",x"49",x"bf",x"f4"),
  1640 => (x"70",x"87",x"da",x"d4"),
  1641 => (x"87",x"c4",x"05",x"98"),
  1642 => (x"4b",x"fe",x"e6",x"c1"),
  1643 => (x"d8",x"ff",x"48",x"73"),
  1644 => (x"52",x"4f",x"87",x"fd"),
  1645 => (x"20",x"20",x"43",x"49"),
  1646 => (x"46",x"43",x"20",x"20"),
  1647 => (x"4f",x"52",x"00",x"47"),
  1648 => (x"6f",x"6c",x"20",x"4d"),
  1649 => (x"6e",x"69",x"64",x"61"),
  1650 => (x"61",x"66",x"20",x"67"),
  1651 => (x"64",x"65",x"6c",x"69"),
  1652 => (x"c6",x"c8",x"1e",x"00"),
  1653 => (x"fd",x"49",x"c1",x"87"),
  1654 => (x"e3",x"fe",x"87",x"ef"),
  1655 => (x"98",x"70",x"87",x"f1"),
  1656 => (x"fe",x"87",x"cd",x"02"),
  1657 => (x"70",x"87",x"ec",x"ec"),
  1658 => (x"87",x"c4",x"02",x"98"),
  1659 => (x"87",x"c2",x"4a",x"c1"),
  1660 => (x"9a",x"72",x"4a",x"c0"),
  1661 => (x"c0",x"87",x"ce",x"05"),
  1662 => (x"e1",x"e8",x"c1",x"1e"),
  1663 => (x"e9",x"f2",x"c0",x"49"),
  1664 => (x"fe",x"86",x"c4",x"87"),
  1665 => (x"c1",x"1e",x"c0",x"87"),
  1666 => (x"c0",x"49",x"ec",x"e8"),
  1667 => (x"c0",x"87",x"db",x"f2"),
  1668 => (x"87",x"f3",x"fd",x"1e"),
  1669 => (x"f2",x"c0",x"49",x"70"),
  1670 => (x"fd",x"c3",x"87",x"d0"),
  1671 => (x"26",x"8e",x"f8",x"87"),
  1672 => (x"20",x"44",x"53",x"4f"),
  1673 => (x"6c",x"69",x"61",x"66"),
  1674 => (x"00",x"2e",x"64",x"65"),
  1675 => (x"74",x"6f",x"6f",x"42"),
  1676 => (x"2e",x"67",x"6e",x"69"),
  1677 => (x"1e",x"00",x"2e",x"2e"),
  1678 => (x"87",x"cd",x"e7",x"c0"),
  1679 => (x"87",x"f9",x"f5",x"c0"),
  1680 => (x"4f",x"26",x"87",x"f6"),
  1681 => (x"e0",x"f4",x"c2",x"1e"),
  1682 => (x"c2",x"78",x"c0",x"48"),
  1683 => (x"c0",x"48",x"c8",x"f4"),
  1684 => (x"87",x"fd",x"fd",x"78"),
  1685 => (x"48",x"c0",x"87",x"e1"),
  1686 => (x"00",x"00",x"4f",x"26"),
  1687 => (x"00",x"00",x"00",x"01"),
  1688 => (x"20",x"20",x"20",x"20"),
  1689 => (x"20",x"20",x"20",x"20"),
  1690 => (x"20",x"20",x"20",x"20"),
  1691 => (x"69",x"78",x"45",x"20"),
  1692 => (x"20",x"20",x"20",x"74"),
  1693 => (x"20",x"20",x"20",x"20"),
  1694 => (x"20",x"20",x"20",x"20"),
  1695 => (x"80",x"00",x"81",x"20"),
  1696 => (x"20",x"20",x"20",x"20"),
  1697 => (x"20",x"20",x"20",x"20"),
  1698 => (x"20",x"20",x"20",x"20"),
  1699 => (x"6b",x"63",x"61",x"42"),
  1700 => (x"00",x"10",x"94",x"00"),
  1701 => (x"00",x"2d",x"34",x"00"),
  1702 => (x"00",x"00",x"00",x"00"),
  1703 => (x"00",x"00",x"10",x"94"),
  1704 => (x"00",x"00",x"2d",x"52"),
  1705 => (x"94",x"00",x"00",x"00"),
  1706 => (x"70",x"00",x"00",x"10"),
  1707 => (x"00",x"00",x"00",x"2d"),
  1708 => (x"10",x"94",x"00",x"00"),
  1709 => (x"2d",x"8e",x"00",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"10",x"94",x"00"),
  1712 => (x"00",x"2d",x"ac",x"00"),
  1713 => (x"00",x"00",x"00",x"00"),
  1714 => (x"00",x"00",x"10",x"94"),
  1715 => (x"00",x"00",x"2d",x"ca"),
  1716 => (x"94",x"00",x"00",x"00"),
  1717 => (x"e8",x"00",x"00",x"10"),
  1718 => (x"00",x"00",x"00",x"2d"),
  1719 => (x"12",x"d3",x"00",x"00"),
  1720 => (x"00",x"00",x"00",x"00"),
  1721 => (x"00",x"00",x"00",x"00"),
  1722 => (x"00",x"13",x"a3",x"00"),
  1723 => (x"00",x"00",x"00",x"00"),
  1724 => (x"00",x"00",x"00",x"00"),
  1725 => (x"00",x"00",x"1a",x"f8"),
  1726 => (x"54",x"4f",x"4f",x"42"),
  1727 => (x"20",x"20",x"20",x"20"),
  1728 => (x"00",x"4d",x"4f",x"52"),
  1729 => (x"48",x"f0",x"fe",x"1e"),
  1730 => (x"09",x"cd",x"78",x"c0"),
  1731 => (x"4f",x"26",x"09",x"79"),
  1732 => (x"f0",x"fe",x"1e",x"1e"),
  1733 => (x"26",x"48",x"7e",x"bf"),
  1734 => (x"fe",x"1e",x"4f",x"26"),
  1735 => (x"78",x"c1",x"48",x"f0"),
  1736 => (x"fe",x"1e",x"4f",x"26"),
  1737 => (x"78",x"c0",x"48",x"f0"),
  1738 => (x"71",x"1e",x"4f",x"26"),
  1739 => (x"52",x"52",x"c0",x"4a"),
  1740 => (x"5e",x"0e",x"4f",x"26"),
  1741 => (x"0e",x"5d",x"5c",x"5b"),
  1742 => (x"4d",x"71",x"86",x"f4"),
  1743 => (x"c1",x"7e",x"6d",x"97"),
  1744 => (x"6c",x"97",x"4c",x"a5"),
  1745 => (x"58",x"a6",x"c8",x"48"),
  1746 => (x"66",x"c4",x"48",x"6e"),
  1747 => (x"87",x"c5",x"05",x"a8"),
  1748 => (x"e6",x"c0",x"48",x"ff"),
  1749 => (x"87",x"ca",x"ff",x"87"),
  1750 => (x"97",x"49",x"a5",x"c2"),
  1751 => (x"a3",x"71",x"4b",x"6c"),
  1752 => (x"4b",x"6b",x"97",x"4b"),
  1753 => (x"6e",x"7e",x"6c",x"97"),
  1754 => (x"c8",x"80",x"c1",x"48"),
  1755 => (x"98",x"c7",x"58",x"a6"),
  1756 => (x"70",x"58",x"a6",x"cc"),
  1757 => (x"e1",x"fe",x"7c",x"97"),
  1758 => (x"f4",x"48",x"73",x"87"),
  1759 => (x"26",x"4d",x"26",x"8e"),
  1760 => (x"26",x"4b",x"26",x"4c"),
  1761 => (x"5b",x"5e",x"0e",x"4f"),
  1762 => (x"86",x"f4",x"0e",x"5c"),
  1763 => (x"66",x"d8",x"4c",x"71"),
  1764 => (x"9a",x"ff",x"c3",x"4a"),
  1765 => (x"97",x"4b",x"a4",x"c2"),
  1766 => (x"a1",x"73",x"49",x"6c"),
  1767 => (x"97",x"51",x"72",x"49"),
  1768 => (x"48",x"6e",x"7e",x"6c"),
  1769 => (x"a6",x"c8",x"80",x"c1"),
  1770 => (x"cc",x"98",x"c7",x"58"),
  1771 => (x"54",x"70",x"58",x"a6"),
  1772 => (x"ca",x"ff",x"8e",x"f4"),
  1773 => (x"fd",x"1e",x"1e",x"87"),
  1774 => (x"bf",x"e0",x"87",x"e8"),
  1775 => (x"e0",x"c0",x"49",x"4a"),
  1776 => (x"cb",x"02",x"99",x"c0"),
  1777 => (x"c2",x"1e",x"72",x"87"),
  1778 => (x"fe",x"49",x"c6",x"f8"),
  1779 => (x"86",x"c4",x"87",x"f7"),
  1780 => (x"70",x"87",x"fd",x"fc"),
  1781 => (x"87",x"c2",x"fd",x"7e"),
  1782 => (x"1e",x"4f",x"26",x"26"),
  1783 => (x"49",x"c6",x"f8",x"c2"),
  1784 => (x"c1",x"87",x"c7",x"fd"),
  1785 => (x"fc",x"49",x"f5",x"ee"),
  1786 => (x"f7",x"c3",x"87",x"da"),
  1787 => (x"0e",x"4f",x"26",x"87"),
  1788 => (x"5d",x"5c",x"5b",x"5e"),
  1789 => (x"c2",x"4d",x"71",x"0e"),
  1790 => (x"fc",x"49",x"c6",x"f8"),
  1791 => (x"4b",x"70",x"87",x"f4"),
  1792 => (x"04",x"ab",x"b7",x"c0"),
  1793 => (x"c3",x"87",x"c2",x"c3"),
  1794 => (x"c9",x"05",x"ab",x"f0"),
  1795 => (x"d3",x"f3",x"c1",x"87"),
  1796 => (x"c2",x"78",x"c1",x"48"),
  1797 => (x"e0",x"c3",x"87",x"e3"),
  1798 => (x"87",x"c9",x"05",x"ab"),
  1799 => (x"48",x"d7",x"f3",x"c1"),
  1800 => (x"d4",x"c2",x"78",x"c1"),
  1801 => (x"d7",x"f3",x"c1",x"87"),
  1802 => (x"87",x"c6",x"02",x"bf"),
  1803 => (x"4c",x"a3",x"c0",x"c2"),
  1804 => (x"4c",x"73",x"87",x"c2"),
  1805 => (x"bf",x"d3",x"f3",x"c1"),
  1806 => (x"87",x"e0",x"c0",x"02"),
  1807 => (x"b7",x"c4",x"49",x"74"),
  1808 => (x"f4",x"c1",x"91",x"29"),
  1809 => (x"4a",x"74",x"81",x"f3"),
  1810 => (x"92",x"c2",x"9a",x"cf"),
  1811 => (x"30",x"72",x"48",x"c1"),
  1812 => (x"ba",x"ff",x"4a",x"70"),
  1813 => (x"98",x"69",x"48",x"72"),
  1814 => (x"87",x"db",x"79",x"70"),
  1815 => (x"b7",x"c4",x"49",x"74"),
  1816 => (x"f4",x"c1",x"91",x"29"),
  1817 => (x"4a",x"74",x"81",x"f3"),
  1818 => (x"92",x"c2",x"9a",x"cf"),
  1819 => (x"30",x"72",x"48",x"c3"),
  1820 => (x"69",x"48",x"4a",x"70"),
  1821 => (x"75",x"79",x"70",x"b0"),
  1822 => (x"f0",x"c0",x"05",x"9d"),
  1823 => (x"48",x"d0",x"ff",x"87"),
  1824 => (x"ff",x"78",x"e1",x"c8"),
  1825 => (x"78",x"c5",x"48",x"d4"),
  1826 => (x"bf",x"d7",x"f3",x"c1"),
  1827 => (x"c3",x"87",x"c3",x"02"),
  1828 => (x"f3",x"c1",x"78",x"e0"),
  1829 => (x"c6",x"02",x"bf",x"d3"),
  1830 => (x"48",x"d4",x"ff",x"87"),
  1831 => (x"ff",x"78",x"f0",x"c3"),
  1832 => (x"78",x"73",x"48",x"d4"),
  1833 => (x"c8",x"48",x"d0",x"ff"),
  1834 => (x"e0",x"c0",x"78",x"e1"),
  1835 => (x"d7",x"f3",x"c1",x"78"),
  1836 => (x"c1",x"78",x"c0",x"48"),
  1837 => (x"c0",x"48",x"d3",x"f3"),
  1838 => (x"c6",x"f8",x"c2",x"78"),
  1839 => (x"87",x"f2",x"f9",x"49"),
  1840 => (x"b7",x"c0",x"4b",x"70"),
  1841 => (x"fe",x"fc",x"03",x"ab"),
  1842 => (x"26",x"48",x"c0",x"87"),
  1843 => (x"26",x"4c",x"26",x"4d"),
  1844 => (x"00",x"4f",x"26",x"4b"),
  1845 => (x"00",x"00",x"00",x"00"),
  1846 => (x"1e",x"00",x"00",x"00"),
  1847 => (x"fc",x"49",x"4a",x"71"),
  1848 => (x"4f",x"26",x"87",x"cd"),
  1849 => (x"72",x"4a",x"c0",x"1e"),
  1850 => (x"c1",x"91",x"c4",x"49"),
  1851 => (x"c0",x"81",x"f3",x"f4"),
  1852 => (x"d0",x"82",x"c1",x"79"),
  1853 => (x"ee",x"04",x"aa",x"b7"),
  1854 => (x"0e",x"4f",x"26",x"87"),
  1855 => (x"5d",x"5c",x"5b",x"5e"),
  1856 => (x"f8",x"4d",x"71",x"0e"),
  1857 => (x"4a",x"75",x"87",x"dc"),
  1858 => (x"92",x"2a",x"b7",x"c4"),
  1859 => (x"82",x"f3",x"f4",x"c1"),
  1860 => (x"9c",x"cf",x"4c",x"75"),
  1861 => (x"49",x"6a",x"94",x"c2"),
  1862 => (x"c3",x"2b",x"74",x"4b"),
  1863 => (x"74",x"48",x"c2",x"9b"),
  1864 => (x"ff",x"4c",x"70",x"30"),
  1865 => (x"71",x"48",x"74",x"bc"),
  1866 => (x"f7",x"7a",x"70",x"98"),
  1867 => (x"48",x"73",x"87",x"ec"),
  1868 => (x"00",x"87",x"d8",x"fe"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"00",x"00"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"00",x"00"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"00",x"00"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"1e",x"00",x"00",x"00"),
  1885 => (x"c8",x"48",x"d0",x"ff"),
  1886 => (x"48",x"71",x"78",x"e1"),
  1887 => (x"78",x"08",x"d4",x"ff"),
  1888 => (x"ff",x"1e",x"4f",x"26"),
  1889 => (x"e1",x"c8",x"48",x"d0"),
  1890 => (x"ff",x"48",x"71",x"78"),
  1891 => (x"c4",x"78",x"08",x"d4"),
  1892 => (x"d4",x"ff",x"48",x"66"),
  1893 => (x"4f",x"26",x"78",x"08"),
  1894 => (x"c4",x"4a",x"71",x"1e"),
  1895 => (x"72",x"1e",x"49",x"66"),
  1896 => (x"87",x"de",x"ff",x"49"),
  1897 => (x"c0",x"48",x"d0",x"ff"),
  1898 => (x"26",x"26",x"78",x"e0"),
  1899 => (x"1e",x"73",x"1e",x"4f"),
  1900 => (x"66",x"c8",x"4b",x"71"),
  1901 => (x"4a",x"73",x"1e",x"49"),
  1902 => (x"49",x"a2",x"e0",x"c1"),
  1903 => (x"26",x"87",x"d9",x"ff"),
  1904 => (x"4d",x"26",x"87",x"c4"),
  1905 => (x"4b",x"26",x"4c",x"26"),
  1906 => (x"73",x"1e",x"4f",x"26"),
  1907 => (x"4b",x"4a",x"71",x"1e"),
  1908 => (x"03",x"ab",x"b7",x"c2"),
  1909 => (x"49",x"a3",x"87",x"c8"),
  1910 => (x"9a",x"ff",x"c3",x"4a"),
  1911 => (x"a3",x"ce",x"87",x"c7"),
  1912 => (x"ff",x"c3",x"4a",x"49"),
  1913 => (x"49",x"66",x"c8",x"9a"),
  1914 => (x"fe",x"49",x"72",x"1e"),
  1915 => (x"ff",x"26",x"87",x"ea"),
  1916 => (x"ff",x"1e",x"87",x"d4"),
  1917 => (x"ff",x"c3",x"4a",x"d4"),
  1918 => (x"48",x"d0",x"ff",x"7a"),
  1919 => (x"de",x"78",x"e1",x"c0"),
  1920 => (x"d0",x"f8",x"c2",x"7a"),
  1921 => (x"48",x"49",x"7a",x"bf"),
  1922 => (x"7a",x"70",x"28",x"c8"),
  1923 => (x"28",x"d0",x"48",x"71"),
  1924 => (x"48",x"71",x"7a",x"70"),
  1925 => (x"7a",x"70",x"28",x"d8"),
  1926 => (x"c0",x"48",x"d0",x"ff"),
  1927 => (x"4f",x"26",x"78",x"e0"),
  1928 => (x"48",x"d0",x"ff",x"1e"),
  1929 => (x"71",x"78",x"c9",x"c8"),
  1930 => (x"08",x"d4",x"ff",x"48"),
  1931 => (x"1e",x"4f",x"26",x"78"),
  1932 => (x"eb",x"49",x"4a",x"71"),
  1933 => (x"48",x"d0",x"ff",x"87"),
  1934 => (x"4f",x"26",x"78",x"c8"),
  1935 => (x"71",x"1e",x"73",x"1e"),
  1936 => (x"e0",x"f8",x"c2",x"4b"),
  1937 => (x"87",x"c3",x"02",x"bf"),
  1938 => (x"ff",x"87",x"eb",x"c2"),
  1939 => (x"c9",x"c8",x"48",x"d0"),
  1940 => (x"c0",x"49",x"73",x"78"),
  1941 => (x"d4",x"ff",x"b1",x"e0"),
  1942 => (x"c2",x"78",x"71",x"48"),
  1943 => (x"c0",x"48",x"d4",x"f8"),
  1944 => (x"02",x"66",x"c8",x"78"),
  1945 => (x"ff",x"c3",x"87",x"c5"),
  1946 => (x"c0",x"87",x"c2",x"49"),
  1947 => (x"dc",x"f8",x"c2",x"49"),
  1948 => (x"02",x"66",x"cc",x"59"),
  1949 => (x"d5",x"c5",x"87",x"c6"),
  1950 => (x"87",x"c4",x"4a",x"d5"),
  1951 => (x"4a",x"ff",x"ff",x"cf"),
  1952 => (x"5a",x"e0",x"f8",x"c2"),
  1953 => (x"48",x"e0",x"f8",x"c2"),
  1954 => (x"87",x"c4",x"78",x"c1"),
  1955 => (x"4c",x"26",x"4d",x"26"),
  1956 => (x"4f",x"26",x"4b",x"26"),
  1957 => (x"5c",x"5b",x"5e",x"0e"),
  1958 => (x"4a",x"71",x"0e",x"5d"),
  1959 => (x"bf",x"dc",x"f8",x"c2"),
  1960 => (x"02",x"9a",x"72",x"4c"),
  1961 => (x"c8",x"49",x"87",x"cb"),
  1962 => (x"f2",x"f8",x"c1",x"91"),
  1963 => (x"c4",x"83",x"71",x"4b"),
  1964 => (x"f2",x"fc",x"c1",x"87"),
  1965 => (x"13",x"4d",x"c0",x"4b"),
  1966 => (x"c2",x"99",x"74",x"49"),
  1967 => (x"b9",x"bf",x"d8",x"f8"),
  1968 => (x"71",x"48",x"d4",x"ff"),
  1969 => (x"2c",x"b7",x"c1",x"78"),
  1970 => (x"ad",x"b7",x"c8",x"85"),
  1971 => (x"c2",x"87",x"e8",x"04"),
  1972 => (x"48",x"bf",x"d4",x"f8"),
  1973 => (x"f8",x"c2",x"80",x"c8"),
  1974 => (x"ef",x"fe",x"58",x"d8"),
  1975 => (x"1e",x"73",x"1e",x"87"),
  1976 => (x"4a",x"13",x"4b",x"71"),
  1977 => (x"87",x"cb",x"02",x"9a"),
  1978 => (x"e7",x"fe",x"49",x"72"),
  1979 => (x"9a",x"4a",x"13",x"87"),
  1980 => (x"fe",x"87",x"f5",x"05"),
  1981 => (x"c2",x"1e",x"87",x"da"),
  1982 => (x"49",x"bf",x"d4",x"f8"),
  1983 => (x"48",x"d4",x"f8",x"c2"),
  1984 => (x"c4",x"78",x"a1",x"c1"),
  1985 => (x"03",x"a9",x"b7",x"c0"),
  1986 => (x"d4",x"ff",x"87",x"db"),
  1987 => (x"d8",x"f8",x"c2",x"48"),
  1988 => (x"f8",x"c2",x"78",x"bf"),
  1989 => (x"c2",x"49",x"bf",x"d4"),
  1990 => (x"c1",x"48",x"d4",x"f8"),
  1991 => (x"c0",x"c4",x"78",x"a1"),
  1992 => (x"e5",x"04",x"a9",x"b7"),
  1993 => (x"48",x"d0",x"ff",x"87"),
  1994 => (x"f8",x"c2",x"78",x"c8"),
  1995 => (x"78",x"c0",x"48",x"e0"),
  1996 => (x"00",x"00",x"4f",x"26"),
  1997 => (x"00",x"00",x"00",x"00"),
  1998 => (x"00",x"00",x"00",x"00"),
  1999 => (x"00",x"5f",x"5f",x"00"),
  2000 => (x"03",x"00",x"00",x"00"),
  2001 => (x"03",x"03",x"00",x"03"),
  2002 => (x"7f",x"14",x"00",x"00"),
  2003 => (x"7f",x"7f",x"14",x"7f"),
  2004 => (x"24",x"00",x"00",x"14"),
  2005 => (x"3a",x"6b",x"6b",x"2e"),
  2006 => (x"6a",x"4c",x"00",x"12"),
  2007 => (x"56",x"6c",x"18",x"36"),
  2008 => (x"7e",x"30",x"00",x"32"),
  2009 => (x"3a",x"77",x"59",x"4f"),
  2010 => (x"00",x"00",x"40",x"68"),
  2011 => (x"00",x"03",x"07",x"04"),
  2012 => (x"00",x"00",x"00",x"00"),
  2013 => (x"41",x"63",x"3e",x"1c"),
  2014 => (x"00",x"00",x"00",x"00"),
  2015 => (x"1c",x"3e",x"63",x"41"),
  2016 => (x"2a",x"08",x"00",x"00"),
  2017 => (x"3e",x"1c",x"1c",x"3e"),
  2018 => (x"08",x"00",x"08",x"2a"),
  2019 => (x"08",x"3e",x"3e",x"08"),
  2020 => (x"00",x"00",x"00",x"08"),
  2021 => (x"00",x"60",x"e0",x"80"),
  2022 => (x"08",x"00",x"00",x"00"),
  2023 => (x"08",x"08",x"08",x"08"),
  2024 => (x"00",x"00",x"00",x"08"),
  2025 => (x"00",x"60",x"60",x"00"),
  2026 => (x"60",x"40",x"00",x"00"),
  2027 => (x"06",x"0c",x"18",x"30"),
  2028 => (x"3e",x"00",x"01",x"03"),
  2029 => (x"7f",x"4d",x"59",x"7f"),
  2030 => (x"04",x"00",x"00",x"3e"),
  2031 => (x"00",x"7f",x"7f",x"06"),
  2032 => (x"42",x"00",x"00",x"00"),
  2033 => (x"4f",x"59",x"71",x"63"),
  2034 => (x"22",x"00",x"00",x"46"),
  2035 => (x"7f",x"49",x"49",x"63"),
  2036 => (x"1c",x"18",x"00",x"36"),
  2037 => (x"7f",x"7f",x"13",x"16"),
  2038 => (x"27",x"00",x"00",x"10"),
  2039 => (x"7d",x"45",x"45",x"67"),
  2040 => (x"3c",x"00",x"00",x"39"),
  2041 => (x"79",x"49",x"4b",x"7e"),
  2042 => (x"01",x"00",x"00",x"30"),
  2043 => (x"0f",x"79",x"71",x"01"),
  2044 => (x"36",x"00",x"00",x"07"),
  2045 => (x"7f",x"49",x"49",x"7f"),
  2046 => (x"06",x"00",x"00",x"36"),
  2047 => (x"3f",x"69",x"49",x"4f"),
  2048 => (x"00",x"00",x"00",x"1e"),
  2049 => (x"00",x"66",x"66",x"00"),
  2050 => (x"00",x"00",x"00",x"00"),
  2051 => (x"00",x"66",x"e6",x"80"),
  2052 => (x"08",x"00",x"00",x"00"),
  2053 => (x"22",x"14",x"14",x"08"),
  2054 => (x"14",x"00",x"00",x"22"),
  2055 => (x"14",x"14",x"14",x"14"),
  2056 => (x"22",x"00",x"00",x"14"),
  2057 => (x"08",x"14",x"14",x"22"),
  2058 => (x"02",x"00",x"00",x"08"),
  2059 => (x"0f",x"59",x"51",x"03"),
  2060 => (x"7f",x"3e",x"00",x"06"),
  2061 => (x"1f",x"55",x"5d",x"41"),
  2062 => (x"7e",x"00",x"00",x"1e"),
  2063 => (x"7f",x"09",x"09",x"7f"),
  2064 => (x"7f",x"00",x"00",x"7e"),
  2065 => (x"7f",x"49",x"49",x"7f"),
  2066 => (x"1c",x"00",x"00",x"36"),
  2067 => (x"41",x"41",x"63",x"3e"),
  2068 => (x"7f",x"00",x"00",x"41"),
  2069 => (x"3e",x"63",x"41",x"7f"),
  2070 => (x"7f",x"00",x"00",x"1c"),
  2071 => (x"41",x"49",x"49",x"7f"),
  2072 => (x"7f",x"00",x"00",x"41"),
  2073 => (x"01",x"09",x"09",x"7f"),
  2074 => (x"3e",x"00",x"00",x"01"),
  2075 => (x"7b",x"49",x"41",x"7f"),
  2076 => (x"7f",x"00",x"00",x"7a"),
  2077 => (x"7f",x"08",x"08",x"7f"),
  2078 => (x"00",x"00",x"00",x"7f"),
  2079 => (x"41",x"7f",x"7f",x"41"),
  2080 => (x"20",x"00",x"00",x"00"),
  2081 => (x"7f",x"40",x"40",x"60"),
  2082 => (x"7f",x"7f",x"00",x"3f"),
  2083 => (x"63",x"36",x"1c",x"08"),
  2084 => (x"7f",x"00",x"00",x"41"),
  2085 => (x"40",x"40",x"40",x"7f"),
  2086 => (x"7f",x"7f",x"00",x"40"),
  2087 => (x"7f",x"06",x"0c",x"06"),
  2088 => (x"7f",x"7f",x"00",x"7f"),
  2089 => (x"7f",x"18",x"0c",x"06"),
  2090 => (x"3e",x"00",x"00",x"7f"),
  2091 => (x"7f",x"41",x"41",x"7f"),
  2092 => (x"7f",x"00",x"00",x"3e"),
  2093 => (x"0f",x"09",x"09",x"7f"),
  2094 => (x"7f",x"3e",x"00",x"06"),
  2095 => (x"7e",x"7f",x"61",x"41"),
  2096 => (x"7f",x"00",x"00",x"40"),
  2097 => (x"7f",x"19",x"09",x"7f"),
  2098 => (x"26",x"00",x"00",x"66"),
  2099 => (x"7b",x"59",x"4d",x"6f"),
  2100 => (x"01",x"00",x"00",x"32"),
  2101 => (x"01",x"7f",x"7f",x"01"),
  2102 => (x"3f",x"00",x"00",x"01"),
  2103 => (x"7f",x"40",x"40",x"7f"),
  2104 => (x"0f",x"00",x"00",x"3f"),
  2105 => (x"3f",x"70",x"70",x"3f"),
  2106 => (x"7f",x"7f",x"00",x"0f"),
  2107 => (x"7f",x"30",x"18",x"30"),
  2108 => (x"63",x"41",x"00",x"7f"),
  2109 => (x"36",x"1c",x"1c",x"36"),
  2110 => (x"03",x"01",x"41",x"63"),
  2111 => (x"06",x"7c",x"7c",x"06"),
  2112 => (x"71",x"61",x"01",x"03"),
  2113 => (x"43",x"47",x"4d",x"59"),
  2114 => (x"00",x"00",x"00",x"41"),
  2115 => (x"41",x"41",x"7f",x"7f"),
  2116 => (x"03",x"01",x"00",x"00"),
  2117 => (x"30",x"18",x"0c",x"06"),
  2118 => (x"00",x"00",x"40",x"60"),
  2119 => (x"7f",x"7f",x"41",x"41"),
  2120 => (x"0c",x"08",x"00",x"00"),
  2121 => (x"0c",x"06",x"03",x"06"),
  2122 => (x"80",x"80",x"00",x"08"),
  2123 => (x"80",x"80",x"80",x"80"),
  2124 => (x"00",x"00",x"00",x"80"),
  2125 => (x"04",x"07",x"03",x"00"),
  2126 => (x"20",x"00",x"00",x"00"),
  2127 => (x"7c",x"54",x"54",x"74"),
  2128 => (x"7f",x"00",x"00",x"78"),
  2129 => (x"7c",x"44",x"44",x"7f"),
  2130 => (x"38",x"00",x"00",x"38"),
  2131 => (x"44",x"44",x"44",x"7c"),
  2132 => (x"38",x"00",x"00",x"00"),
  2133 => (x"7f",x"44",x"44",x"7c"),
  2134 => (x"38",x"00",x"00",x"7f"),
  2135 => (x"5c",x"54",x"54",x"7c"),
  2136 => (x"04",x"00",x"00",x"18"),
  2137 => (x"05",x"05",x"7f",x"7e"),
  2138 => (x"18",x"00",x"00",x"00"),
  2139 => (x"fc",x"a4",x"a4",x"bc"),
  2140 => (x"7f",x"00",x"00",x"7c"),
  2141 => (x"7c",x"04",x"04",x"7f"),
  2142 => (x"00",x"00",x"00",x"78"),
  2143 => (x"40",x"7d",x"3d",x"00"),
  2144 => (x"80",x"00",x"00",x"00"),
  2145 => (x"7d",x"fd",x"80",x"80"),
  2146 => (x"7f",x"00",x"00",x"00"),
  2147 => (x"6c",x"38",x"10",x"7f"),
  2148 => (x"00",x"00",x"00",x"44"),
  2149 => (x"40",x"7f",x"3f",x"00"),
  2150 => (x"7c",x"7c",x"00",x"00"),
  2151 => (x"7c",x"0c",x"18",x"0c"),
  2152 => (x"7c",x"00",x"00",x"78"),
  2153 => (x"7c",x"04",x"04",x"7c"),
  2154 => (x"38",x"00",x"00",x"78"),
  2155 => (x"7c",x"44",x"44",x"7c"),
  2156 => (x"fc",x"00",x"00",x"38"),
  2157 => (x"3c",x"24",x"24",x"fc"),
  2158 => (x"18",x"00",x"00",x"18"),
  2159 => (x"fc",x"24",x"24",x"3c"),
  2160 => (x"7c",x"00",x"00",x"fc"),
  2161 => (x"0c",x"04",x"04",x"7c"),
  2162 => (x"48",x"00",x"00",x"08"),
  2163 => (x"74",x"54",x"54",x"5c"),
  2164 => (x"04",x"00",x"00",x"20"),
  2165 => (x"44",x"44",x"7f",x"3f"),
  2166 => (x"3c",x"00",x"00",x"00"),
  2167 => (x"7c",x"40",x"40",x"7c"),
  2168 => (x"1c",x"00",x"00",x"7c"),
  2169 => (x"3c",x"60",x"60",x"3c"),
  2170 => (x"7c",x"3c",x"00",x"1c"),
  2171 => (x"7c",x"60",x"30",x"60"),
  2172 => (x"6c",x"44",x"00",x"3c"),
  2173 => (x"6c",x"38",x"10",x"38"),
  2174 => (x"1c",x"00",x"00",x"44"),
  2175 => (x"3c",x"60",x"e0",x"bc"),
  2176 => (x"44",x"00",x"00",x"1c"),
  2177 => (x"4c",x"5c",x"74",x"64"),
  2178 => (x"08",x"00",x"00",x"44"),
  2179 => (x"41",x"77",x"3e",x"08"),
  2180 => (x"00",x"00",x"00",x"41"),
  2181 => (x"00",x"7f",x"7f",x"00"),
  2182 => (x"41",x"00",x"00",x"00"),
  2183 => (x"08",x"3e",x"77",x"41"),
  2184 => (x"01",x"02",x"00",x"08"),
  2185 => (x"02",x"02",x"03",x"01"),
  2186 => (x"7f",x"7f",x"00",x"01"),
  2187 => (x"7f",x"7f",x"7f",x"7f"),
  2188 => (x"08",x"08",x"00",x"7f"),
  2189 => (x"3e",x"3e",x"1c",x"1c"),
  2190 => (x"7f",x"7f",x"7f",x"7f"),
  2191 => (x"1c",x"1c",x"3e",x"3e"),
  2192 => (x"10",x"00",x"08",x"08"),
  2193 => (x"18",x"7c",x"7c",x"18"),
  2194 => (x"10",x"00",x"00",x"10"),
  2195 => (x"30",x"7c",x"7c",x"30"),
  2196 => (x"30",x"10",x"00",x"10"),
  2197 => (x"1e",x"78",x"60",x"60"),
  2198 => (x"66",x"42",x"00",x"06"),
  2199 => (x"66",x"3c",x"18",x"3c"),
  2200 => (x"38",x"78",x"00",x"42"),
  2201 => (x"6c",x"c6",x"c2",x"6a"),
  2202 => (x"00",x"60",x"00",x"38"),
  2203 => (x"00",x"00",x"60",x"00"),
  2204 => (x"5e",x"0e",x"00",x"60"),
  2205 => (x"0e",x"5d",x"5c",x"5b"),
  2206 => (x"c2",x"4c",x"71",x"1e"),
  2207 => (x"4d",x"bf",x"f1",x"f8"),
  2208 => (x"1e",x"c0",x"4b",x"c0"),
  2209 => (x"c7",x"02",x"ab",x"74"),
  2210 => (x"48",x"a6",x"c4",x"87"),
  2211 => (x"87",x"c5",x"78",x"c0"),
  2212 => (x"c1",x"48",x"a6",x"c4"),
  2213 => (x"1e",x"66",x"c4",x"78"),
  2214 => (x"df",x"ee",x"49",x"73"),
  2215 => (x"c0",x"86",x"c8",x"87"),
  2216 => (x"ef",x"ef",x"49",x"e0"),
  2217 => (x"4a",x"a5",x"c4",x"87"),
  2218 => (x"f0",x"f0",x"49",x"6a"),
  2219 => (x"87",x"c6",x"f1",x"87"),
  2220 => (x"83",x"c1",x"85",x"cb"),
  2221 => (x"04",x"ab",x"b7",x"c8"),
  2222 => (x"26",x"87",x"c7",x"ff"),
  2223 => (x"4c",x"26",x"4d",x"26"),
  2224 => (x"4f",x"26",x"4b",x"26"),
  2225 => (x"c2",x"4a",x"71",x"1e"),
  2226 => (x"c2",x"5a",x"f5",x"f8"),
  2227 => (x"c7",x"48",x"f5",x"f8"),
  2228 => (x"dd",x"fe",x"49",x"78"),
  2229 => (x"1e",x"4f",x"26",x"87"),
  2230 => (x"4a",x"71",x"1e",x"73"),
  2231 => (x"03",x"aa",x"b7",x"c0"),
  2232 => (x"dc",x"c2",x"87",x"d3"),
  2233 => (x"c4",x"05",x"bf",x"d8"),
  2234 => (x"c2",x"4b",x"c1",x"87"),
  2235 => (x"c2",x"4b",x"c0",x"87"),
  2236 => (x"c4",x"5b",x"dc",x"dc"),
  2237 => (x"dc",x"dc",x"c2",x"87"),
  2238 => (x"d8",x"dc",x"c2",x"5a"),
  2239 => (x"9a",x"c1",x"4a",x"bf"),
  2240 => (x"49",x"a2",x"c0",x"c1"),
  2241 => (x"c2",x"87",x"e8",x"ec"),
  2242 => (x"49",x"bf",x"c0",x"dc"),
  2243 => (x"bf",x"d8",x"dc",x"c2"),
  2244 => (x"71",x"48",x"fc",x"b1"),
  2245 => (x"87",x"e8",x"fe",x"78"),
  2246 => (x"c4",x"4a",x"71",x"1e"),
  2247 => (x"49",x"72",x"1e",x"66"),
  2248 => (x"26",x"87",x"e7",x"ea"),
  2249 => (x"71",x"1e",x"4f",x"26"),
  2250 => (x"48",x"d4",x"ff",x"4a"),
  2251 => (x"ff",x"78",x"ff",x"c3"),
  2252 => (x"e1",x"c0",x"48",x"d0"),
  2253 => (x"48",x"d4",x"ff",x"78"),
  2254 => (x"49",x"72",x"78",x"c1"),
  2255 => (x"78",x"71",x"31",x"c4"),
  2256 => (x"c0",x"48",x"d0",x"ff"),
  2257 => (x"4f",x"26",x"78",x"e0"),
  2258 => (x"d8",x"dc",x"c2",x"1e"),
  2259 => (x"ca",x"e6",x"49",x"bf"),
  2260 => (x"e9",x"f8",x"c2",x"87"),
  2261 => (x"78",x"bf",x"e8",x"48"),
  2262 => (x"48",x"e5",x"f8",x"c2"),
  2263 => (x"c2",x"78",x"bf",x"ec"),
  2264 => (x"4a",x"bf",x"e9",x"f8"),
  2265 => (x"99",x"ff",x"c3",x"49"),
  2266 => (x"72",x"2a",x"b7",x"c8"),
  2267 => (x"c2",x"b0",x"71",x"48"),
  2268 => (x"26",x"58",x"f1",x"f8"),
  2269 => (x"5b",x"5e",x"0e",x"4f"),
  2270 => (x"71",x"0e",x"5d",x"5c"),
  2271 => (x"87",x"c8",x"ff",x"4b"),
  2272 => (x"48",x"e4",x"f8",x"c2"),
  2273 => (x"49",x"73",x"50",x"c0"),
  2274 => (x"70",x"87",x"f0",x"e5"),
  2275 => (x"9c",x"c2",x"4c",x"49"),
  2276 => (x"ce",x"49",x"ee",x"cb"),
  2277 => (x"49",x"70",x"87",x"ca"),
  2278 => (x"e4",x"f8",x"c2",x"4d"),
  2279 => (x"c1",x"05",x"bf",x"97"),
  2280 => (x"66",x"d0",x"87",x"e2"),
  2281 => (x"ed",x"f8",x"c2",x"49"),
  2282 => (x"d6",x"05",x"99",x"bf"),
  2283 => (x"49",x"66",x"d4",x"87"),
  2284 => (x"bf",x"e5",x"f8",x"c2"),
  2285 => (x"87",x"cb",x"05",x"99"),
  2286 => (x"fe",x"e4",x"49",x"73"),
  2287 => (x"02",x"98",x"70",x"87"),
  2288 => (x"c1",x"87",x"c1",x"c1"),
  2289 => (x"87",x"c0",x"fe",x"4c"),
  2290 => (x"df",x"cd",x"49",x"75"),
  2291 => (x"02",x"98",x"70",x"87"),
  2292 => (x"f8",x"c2",x"87",x"c6"),
  2293 => (x"50",x"c1",x"48",x"e4"),
  2294 => (x"97",x"e4",x"f8",x"c2"),
  2295 => (x"e3",x"c0",x"05",x"bf"),
  2296 => (x"ed",x"f8",x"c2",x"87"),
  2297 => (x"66",x"d0",x"49",x"bf"),
  2298 => (x"d6",x"ff",x"05",x"99"),
  2299 => (x"e5",x"f8",x"c2",x"87"),
  2300 => (x"66",x"d4",x"49",x"bf"),
  2301 => (x"ca",x"ff",x"05",x"99"),
  2302 => (x"e3",x"49",x"73",x"87"),
  2303 => (x"98",x"70",x"87",x"fd"),
  2304 => (x"87",x"ff",x"fe",x"05"),
  2305 => (x"f3",x"fa",x"48",x"74"),
  2306 => (x"5b",x"5e",x"0e",x"87"),
  2307 => (x"f4",x"0e",x"5d",x"5c"),
  2308 => (x"4c",x"4d",x"c0",x"86"),
  2309 => (x"c4",x"7e",x"bf",x"ec"),
  2310 => (x"f8",x"c2",x"48",x"a6"),
  2311 => (x"c0",x"78",x"bf",x"f1"),
  2312 => (x"f7",x"c1",x"1e",x"1e"),
  2313 => (x"87",x"cd",x"fd",x"49"),
  2314 => (x"98",x"70",x"86",x"c8"),
  2315 => (x"87",x"f3",x"c0",x"02"),
  2316 => (x"bf",x"c0",x"dc",x"c2"),
  2317 => (x"c1",x"87",x"c4",x"05"),
  2318 => (x"c0",x"87",x"c2",x"7e"),
  2319 => (x"c0",x"dc",x"c2",x"7e"),
  2320 => (x"ca",x"78",x"6e",x"48"),
  2321 => (x"66",x"c4",x"1e",x"fc"),
  2322 => (x"c4",x"87",x"c9",x"02"),
  2323 => (x"da",x"c2",x"48",x"a6"),
  2324 => (x"87",x"c7",x"78",x"d3"),
  2325 => (x"c2",x"48",x"a6",x"c4"),
  2326 => (x"c4",x"78",x"de",x"da"),
  2327 => (x"c9",x"c9",x"49",x"66"),
  2328 => (x"c1",x"86",x"c4",x"87"),
  2329 => (x"c7",x"1e",x"c0",x"1e"),
  2330 => (x"87",x"c9",x"fc",x"49"),
  2331 => (x"98",x"70",x"86",x"c8"),
  2332 => (x"ff",x"87",x"cd",x"02"),
  2333 => (x"87",x"df",x"f9",x"49"),
  2334 => (x"e1",x"49",x"da",x"c1"),
  2335 => (x"4d",x"c1",x"87",x"fd"),
  2336 => (x"97",x"e4",x"f8",x"c2"),
  2337 => (x"87",x"cf",x"02",x"bf"),
  2338 => (x"bf",x"fc",x"db",x"c2"),
  2339 => (x"c2",x"b9",x"c1",x"49"),
  2340 => (x"71",x"59",x"c0",x"dc"),
  2341 => (x"c2",x"87",x"cf",x"fa"),
  2342 => (x"4b",x"bf",x"e9",x"f8"),
  2343 => (x"bf",x"d8",x"dc",x"c2"),
  2344 => (x"87",x"e1",x"c1",x"05"),
  2345 => (x"bf",x"c0",x"dc",x"c2"),
  2346 => (x"87",x"f0",x"c0",x"02"),
  2347 => (x"c8",x"48",x"a6",x"c4"),
  2348 => (x"c2",x"78",x"c0",x"c0"),
  2349 => (x"6e",x"7e",x"c4",x"dc"),
  2350 => (x"6e",x"49",x"bf",x"97"),
  2351 => (x"70",x"80",x"c1",x"48"),
  2352 => (x"f6",x"e0",x"71",x"7e"),
  2353 => (x"02",x"98",x"70",x"87"),
  2354 => (x"66",x"c4",x"87",x"c3"),
  2355 => (x"48",x"66",x"c4",x"b3"),
  2356 => (x"c8",x"28",x"b7",x"c1"),
  2357 => (x"98",x"70",x"58",x"a6"),
  2358 => (x"87",x"db",x"ff",x"05"),
  2359 => (x"e0",x"49",x"fd",x"c3"),
  2360 => (x"fa",x"c3",x"87",x"d9"),
  2361 => (x"87",x"d3",x"e0",x"49"),
  2362 => (x"ff",x"c3",x"49",x"73"),
  2363 => (x"c0",x"1e",x"71",x"99"),
  2364 => (x"87",x"e4",x"f8",x"49"),
  2365 => (x"b7",x"c8",x"49",x"73"),
  2366 => (x"c1",x"1e",x"71",x"29"),
  2367 => (x"87",x"d8",x"f8",x"49"),
  2368 => (x"c9",x"c6",x"86",x"c8"),
  2369 => (x"ed",x"f8",x"c2",x"87"),
  2370 => (x"02",x"9b",x"4b",x"bf"),
  2371 => (x"dc",x"c2",x"87",x"df"),
  2372 => (x"c8",x"49",x"bf",x"d4"),
  2373 => (x"98",x"70",x"87",x"d6"),
  2374 => (x"87",x"c4",x"c0",x"05"),
  2375 => (x"87",x"d3",x"4b",x"c0"),
  2376 => (x"c7",x"49",x"e0",x"c2"),
  2377 => (x"dc",x"c2",x"87",x"fa"),
  2378 => (x"c6",x"c0",x"58",x"d8"),
  2379 => (x"d4",x"dc",x"c2",x"87"),
  2380 => (x"73",x"78",x"c0",x"48"),
  2381 => (x"05",x"99",x"c2",x"49"),
  2382 => (x"c3",x"87",x"cf",x"c0"),
  2383 => (x"de",x"ff",x"49",x"eb"),
  2384 => (x"49",x"70",x"87",x"f9"),
  2385 => (x"c0",x"02",x"99",x"c2"),
  2386 => (x"4c",x"fb",x"87",x"c2"),
  2387 => (x"99",x"c1",x"49",x"73"),
  2388 => (x"87",x"cf",x"c0",x"05"),
  2389 => (x"ff",x"49",x"f4",x"c3"),
  2390 => (x"70",x"87",x"e0",x"de"),
  2391 => (x"02",x"99",x"c2",x"49"),
  2392 => (x"fa",x"87",x"c2",x"c0"),
  2393 => (x"c8",x"49",x"73",x"4c"),
  2394 => (x"cf",x"c0",x"05",x"99"),
  2395 => (x"49",x"f5",x"c3",x"87"),
  2396 => (x"87",x"c7",x"de",x"ff"),
  2397 => (x"99",x"c2",x"49",x"70"),
  2398 => (x"87",x"d6",x"c0",x"02"),
  2399 => (x"bf",x"f5",x"f8",x"c2"),
  2400 => (x"87",x"ca",x"c0",x"02"),
  2401 => (x"c2",x"88",x"c1",x"48"),
  2402 => (x"c0",x"58",x"f9",x"f8"),
  2403 => (x"4c",x"ff",x"87",x"c2"),
  2404 => (x"49",x"73",x"4d",x"c1"),
  2405 => (x"c0",x"05",x"99",x"c4"),
  2406 => (x"f2",x"c3",x"87",x"cf"),
  2407 => (x"da",x"dd",x"ff",x"49"),
  2408 => (x"c2",x"49",x"70",x"87"),
  2409 => (x"dc",x"c0",x"02",x"99"),
  2410 => (x"f5",x"f8",x"c2",x"87"),
  2411 => (x"c7",x"48",x"7e",x"bf"),
  2412 => (x"c0",x"03",x"a8",x"b7"),
  2413 => (x"48",x"6e",x"87",x"cb"),
  2414 => (x"f8",x"c2",x"80",x"c1"),
  2415 => (x"c2",x"c0",x"58",x"f9"),
  2416 => (x"c1",x"4c",x"fe",x"87"),
  2417 => (x"49",x"fd",x"c3",x"4d"),
  2418 => (x"87",x"ef",x"dc",x"ff"),
  2419 => (x"99",x"c2",x"49",x"70"),
  2420 => (x"87",x"d5",x"c0",x"02"),
  2421 => (x"bf",x"f5",x"f8",x"c2"),
  2422 => (x"87",x"c9",x"c0",x"02"),
  2423 => (x"48",x"f5",x"f8",x"c2"),
  2424 => (x"c2",x"c0",x"78",x"c0"),
  2425 => (x"c1",x"4c",x"fd",x"87"),
  2426 => (x"49",x"fa",x"c3",x"4d"),
  2427 => (x"87",x"cb",x"dc",x"ff"),
  2428 => (x"99",x"c2",x"49",x"70"),
  2429 => (x"87",x"d9",x"c0",x"02"),
  2430 => (x"bf",x"f5",x"f8",x"c2"),
  2431 => (x"a8",x"b7",x"c7",x"48"),
  2432 => (x"87",x"c9",x"c0",x"03"),
  2433 => (x"48",x"f5",x"f8",x"c2"),
  2434 => (x"c2",x"c0",x"78",x"c7"),
  2435 => (x"c1",x"4c",x"fc",x"87"),
  2436 => (x"ac",x"b7",x"c0",x"4d"),
  2437 => (x"87",x"d0",x"c0",x"03"),
  2438 => (x"c1",x"4a",x"66",x"c4"),
  2439 => (x"02",x"6a",x"82",x"d8"),
  2440 => (x"4b",x"87",x"c5",x"c0"),
  2441 => (x"0f",x"73",x"49",x"74"),
  2442 => (x"f0",x"c3",x"1e",x"c0"),
  2443 => (x"49",x"da",x"c1",x"1e"),
  2444 => (x"c8",x"87",x"c2",x"f5"),
  2445 => (x"02",x"98",x"70",x"86"),
  2446 => (x"c8",x"87",x"e0",x"c0"),
  2447 => (x"f8",x"c2",x"48",x"a6"),
  2448 => (x"c8",x"78",x"bf",x"f5"),
  2449 => (x"91",x"cb",x"49",x"66"),
  2450 => (x"71",x"48",x"66",x"c4"),
  2451 => (x"6e",x"7e",x"70",x"80"),
  2452 => (x"c6",x"c0",x"02",x"bf"),
  2453 => (x"66",x"c8",x"4b",x"87"),
  2454 => (x"75",x"0f",x"73",x"49"),
  2455 => (x"c8",x"c0",x"02",x"9d"),
  2456 => (x"f5",x"f8",x"c2",x"87"),
  2457 => (x"c9",x"f0",x"49",x"bf"),
  2458 => (x"dc",x"dc",x"c2",x"87"),
  2459 => (x"dd",x"c0",x"02",x"bf"),
  2460 => (x"f7",x"c2",x"49",x"87"),
  2461 => (x"02",x"98",x"70",x"87"),
  2462 => (x"c2",x"87",x"d3",x"c0"),
  2463 => (x"49",x"bf",x"f5",x"f8"),
  2464 => (x"c0",x"87",x"ef",x"ef"),
  2465 => (x"87",x"cf",x"f1",x"49"),
  2466 => (x"48",x"dc",x"dc",x"c2"),
  2467 => (x"8e",x"f4",x"78",x"c0"),
  2468 => (x"4a",x"87",x"e9",x"f0"),
  2469 => (x"65",x"6b",x"79",x"6f"),
  2470 => (x"6f",x"20",x"73",x"79"),
  2471 => (x"6f",x"4a",x"00",x"6e"),
  2472 => (x"79",x"65",x"6b",x"79"),
  2473 => (x"66",x"6f",x"20",x"73"),
  2474 => (x"5e",x"0e",x"00",x"66"),
  2475 => (x"0e",x"5d",x"5c",x"5b"),
  2476 => (x"c2",x"4c",x"71",x"1e"),
  2477 => (x"49",x"bf",x"f1",x"f8"),
  2478 => (x"4d",x"a1",x"cd",x"c1"),
  2479 => (x"69",x"81",x"d1",x"c1"),
  2480 => (x"02",x"9c",x"74",x"7e"),
  2481 => (x"a5",x"c4",x"87",x"cf"),
  2482 => (x"c2",x"7b",x"74",x"4b"),
  2483 => (x"49",x"bf",x"f1",x"f8"),
  2484 => (x"6e",x"87",x"f1",x"ef"),
  2485 => (x"05",x"9c",x"74",x"7b"),
  2486 => (x"4b",x"c0",x"87",x"c4"),
  2487 => (x"4b",x"c1",x"87",x"c2"),
  2488 => (x"f2",x"ef",x"49",x"73"),
  2489 => (x"02",x"66",x"d4",x"87"),
  2490 => (x"c0",x"49",x"87",x"c8"),
  2491 => (x"4a",x"70",x"87",x"f2"),
  2492 => (x"4a",x"c0",x"87",x"c2"),
  2493 => (x"5a",x"e0",x"dc",x"c2"),
  2494 => (x"87",x"c0",x"ef",x"26"),
  2495 => (x"00",x"00",x"00",x"00"),
  2496 => (x"00",x"00",x"00",x"00"),
  2497 => (x"14",x"11",x"12",x"58"),
  2498 => (x"23",x"1c",x"1b",x"1d"),
  2499 => (x"94",x"91",x"59",x"5a"),
  2500 => (x"f4",x"eb",x"f2",x"f5"),
  2501 => (x"00",x"00",x"00",x"00"),
  2502 => (x"00",x"00",x"00",x"00"),
  2503 => (x"00",x"00",x"00",x"00"),
  2504 => (x"ff",x"4a",x"71",x"1e"),
  2505 => (x"72",x"49",x"bf",x"c8"),
  2506 => (x"4f",x"26",x"48",x"a1"),
  2507 => (x"bf",x"c8",x"ff",x"1e"),
  2508 => (x"c0",x"c0",x"fe",x"89"),
  2509 => (x"a9",x"c0",x"c0",x"c0"),
  2510 => (x"c0",x"87",x"c4",x"01"),
  2511 => (x"c1",x"87",x"c2",x"4a"),
  2512 => (x"26",x"48",x"72",x"4a"),
  2513 => (x"5b",x"5e",x"0e",x"4f"),
  2514 => (x"71",x"0e",x"5d",x"5c"),
  2515 => (x"4c",x"d4",x"ff",x"4b"),
  2516 => (x"c0",x"48",x"66",x"d0"),
  2517 => (x"ff",x"49",x"d6",x"78"),
  2518 => (x"c3",x"87",x"d8",x"d8"),
  2519 => (x"49",x"6c",x"7c",x"ff"),
  2520 => (x"71",x"99",x"ff",x"c3"),
  2521 => (x"f0",x"c3",x"49",x"4d"),
  2522 => (x"a9",x"e0",x"c1",x"99"),
  2523 => (x"c3",x"87",x"cb",x"05"),
  2524 => (x"48",x"6c",x"7c",x"ff"),
  2525 => (x"66",x"d0",x"98",x"c3"),
  2526 => (x"ff",x"c3",x"78",x"08"),
  2527 => (x"49",x"4a",x"6c",x"7c"),
  2528 => (x"ff",x"c3",x"31",x"c8"),
  2529 => (x"71",x"4a",x"6c",x"7c"),
  2530 => (x"c8",x"49",x"72",x"b2"),
  2531 => (x"7c",x"ff",x"c3",x"31"),
  2532 => (x"b2",x"71",x"4a",x"6c"),
  2533 => (x"31",x"c8",x"49",x"72"),
  2534 => (x"6c",x"7c",x"ff",x"c3"),
  2535 => (x"ff",x"b2",x"71",x"4a"),
  2536 => (x"e0",x"c0",x"48",x"d0"),
  2537 => (x"02",x"9b",x"73",x"78"),
  2538 => (x"7b",x"72",x"87",x"c2"),
  2539 => (x"4d",x"26",x"48",x"75"),
  2540 => (x"4b",x"26",x"4c",x"26"),
  2541 => (x"26",x"1e",x"4f",x"26"),
  2542 => (x"5b",x"5e",x"0e",x"4f"),
  2543 => (x"86",x"f8",x"0e",x"5c"),
  2544 => (x"a6",x"c8",x"1e",x"76"),
  2545 => (x"87",x"fd",x"fd",x"49"),
  2546 => (x"4b",x"70",x"86",x"c4"),
  2547 => (x"a8",x"c2",x"48",x"6e"),
  2548 => (x"87",x"f0",x"c2",x"03"),
  2549 => (x"f0",x"c3",x"4a",x"73"),
  2550 => (x"aa",x"d0",x"c1",x"9a"),
  2551 => (x"c1",x"87",x"c7",x"02"),
  2552 => (x"c2",x"05",x"aa",x"e0"),
  2553 => (x"49",x"73",x"87",x"de"),
  2554 => (x"c3",x"02",x"99",x"c8"),
  2555 => (x"87",x"c6",x"ff",x"87"),
  2556 => (x"9c",x"c3",x"4c",x"73"),
  2557 => (x"c1",x"05",x"ac",x"c2"),
  2558 => (x"66",x"c4",x"87",x"c2"),
  2559 => (x"71",x"31",x"c9",x"49"),
  2560 => (x"4a",x"66",x"c4",x"1e"),
  2561 => (x"f8",x"c2",x"92",x"d4"),
  2562 => (x"81",x"72",x"49",x"f9"),
  2563 => (x"87",x"c2",x"c7",x"fe"),
  2564 => (x"d5",x"ff",x"49",x"d8"),
  2565 => (x"c0",x"c8",x"87",x"dd"),
  2566 => (x"d6",x"e7",x"c2",x"1e"),
  2567 => (x"fd",x"e2",x"fd",x"49"),
  2568 => (x"48",x"d0",x"ff",x"87"),
  2569 => (x"c2",x"78",x"e0",x"c0"),
  2570 => (x"cc",x"1e",x"d6",x"e7"),
  2571 => (x"92",x"d4",x"4a",x"66"),
  2572 => (x"49",x"f9",x"f8",x"c2"),
  2573 => (x"c5",x"fe",x"81",x"72"),
  2574 => (x"86",x"cc",x"87",x"c9"),
  2575 => (x"c1",x"05",x"ac",x"c1"),
  2576 => (x"66",x"c4",x"87",x"c2"),
  2577 => (x"71",x"31",x"c9",x"49"),
  2578 => (x"4a",x"66",x"c4",x"1e"),
  2579 => (x"f8",x"c2",x"92",x"d4"),
  2580 => (x"81",x"72",x"49",x"f9"),
  2581 => (x"87",x"fa",x"c5",x"fe"),
  2582 => (x"1e",x"d6",x"e7",x"c2"),
  2583 => (x"d4",x"4a",x"66",x"c8"),
  2584 => (x"f9",x"f8",x"c2",x"92"),
  2585 => (x"fe",x"81",x"72",x"49"),
  2586 => (x"d7",x"87",x"c9",x"c3"),
  2587 => (x"c2",x"d4",x"ff",x"49"),
  2588 => (x"1e",x"c0",x"c8",x"87"),
  2589 => (x"49",x"d6",x"e7",x"c2"),
  2590 => (x"87",x"fb",x"e0",x"fd"),
  2591 => (x"d0",x"ff",x"86",x"cc"),
  2592 => (x"78",x"e0",x"c0",x"48"),
  2593 => (x"e7",x"fc",x"8e",x"f8"),
  2594 => (x"5b",x"5e",x"0e",x"87"),
  2595 => (x"1e",x"0e",x"5d",x"5c"),
  2596 => (x"d4",x"ff",x"4d",x"71"),
  2597 => (x"7e",x"66",x"d4",x"4c"),
  2598 => (x"a8",x"b7",x"c3",x"48"),
  2599 => (x"c0",x"87",x"c5",x"06"),
  2600 => (x"87",x"e2",x"c1",x"48"),
  2601 => (x"d3",x"fe",x"49",x"75"),
  2602 => (x"1e",x"75",x"87",x"f5"),
  2603 => (x"d4",x"4b",x"66",x"c4"),
  2604 => (x"f9",x"f8",x"c2",x"93"),
  2605 => (x"fd",x"49",x"73",x"83"),
  2606 => (x"c8",x"87",x"c5",x"fd"),
  2607 => (x"ff",x"4b",x"6b",x"83"),
  2608 => (x"e1",x"c8",x"48",x"d0"),
  2609 => (x"73",x"7c",x"dd",x"78"),
  2610 => (x"99",x"ff",x"c3",x"49"),
  2611 => (x"49",x"73",x"7c",x"71"),
  2612 => (x"c3",x"29",x"b7",x"c8"),
  2613 => (x"7c",x"71",x"99",x"ff"),
  2614 => (x"b7",x"d0",x"49",x"73"),
  2615 => (x"99",x"ff",x"c3",x"29"),
  2616 => (x"49",x"73",x"7c",x"71"),
  2617 => (x"71",x"29",x"b7",x"d8"),
  2618 => (x"7c",x"7c",x"c0",x"7c"),
  2619 => (x"7c",x"7c",x"7c",x"7c"),
  2620 => (x"7c",x"7c",x"7c",x"7c"),
  2621 => (x"e0",x"c0",x"7c",x"7c"),
  2622 => (x"1e",x"66",x"c4",x"78"),
  2623 => (x"d2",x"ff",x"49",x"dc"),
  2624 => (x"86",x"c8",x"87",x"d6"),
  2625 => (x"fa",x"26",x"48",x"73"),
  2626 => (x"71",x"1e",x"87",x"e4"),
  2627 => (x"49",x"a2",x"c4",x"4a"),
  2628 => (x"48",x"d0",x"f8",x"c2"),
  2629 => (x"db",x"c2",x"78",x"6a"),
  2630 => (x"78",x"69",x"48",x"fc"),
  2631 => (x"bf",x"fc",x"db",x"c2"),
  2632 => (x"87",x"c2",x"e8",x"49"),
  2633 => (x"87",x"ca",x"d3",x"ff"),
  2634 => (x"4f",x"26",x"48",x"c1"),
  2635 => (x"c4",x"4a",x"71",x"1e"),
  2636 => (x"f8",x"c2",x"49",x"a2"),
  2637 => (x"c2",x"7a",x"bf",x"d0"),
  2638 => (x"79",x"bf",x"fc",x"db"),
  2639 => (x"71",x"1e",x"4f",x"26"),
  2640 => (x"c0",x"02",x"9a",x"4a"),
  2641 => (x"c2",x"1e",x"87",x"ec"),
  2642 => (x"fd",x"49",x"cc",x"f4"),
  2643 => (x"c4",x"87",x"f1",x"fa"),
  2644 => (x"02",x"98",x"70",x"86"),
  2645 => (x"e7",x"c2",x"87",x"dc"),
  2646 => (x"f4",x"c2",x"1e",x"d6"),
  2647 => (x"ff",x"fd",x"49",x"cc"),
  2648 => (x"86",x"c4",x"87",x"d2"),
  2649 => (x"c9",x"02",x"98",x"70"),
  2650 => (x"d6",x"e7",x"c2",x"87"),
  2651 => (x"87",x"da",x"fe",x"49"),
  2652 => (x"48",x"c0",x"87",x"c2"),
  2653 => (x"71",x"1e",x"4f",x"26"),
  2654 => (x"c0",x"02",x"9a",x"4a"),
  2655 => (x"c2",x"1e",x"87",x"ee"),
  2656 => (x"fd",x"49",x"cc",x"f4"),
  2657 => (x"c4",x"87",x"f9",x"f9"),
  2658 => (x"02",x"98",x"70",x"86"),
  2659 => (x"e7",x"c2",x"87",x"de"),
  2660 => (x"d7",x"fe",x"49",x"d6"),
  2661 => (x"d6",x"e7",x"c2",x"87"),
  2662 => (x"cc",x"f4",x"c2",x"1e"),
  2663 => (x"e2",x"ff",x"fd",x"49"),
  2664 => (x"70",x"86",x"c4",x"87"),
  2665 => (x"87",x"c4",x"02",x"98"),
  2666 => (x"87",x"c2",x"48",x"c1"),
  2667 => (x"4f",x"26",x"48",x"c0"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

