
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e8",x"c0",x"c3",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"e8",x"c0",x"c3"),
    18 => (x"48",x"c0",x"e8",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"ff",x"e7",x"c2",x"87"),
    25 => (x"fb",x"e7",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"ee",x"c1",x"87",x"f7"),
    29 => (x"e7",x"c2",x"87",x"d1"),
    30 => (x"e7",x"c2",x"4d",x"ff"),
    31 => (x"ad",x"74",x"4c",x"ff"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"86",x"f0",x"0e",x"5d"),
    37 => (x"a6",x"c4",x"4c",x"c0"),
    38 => (x"c0",x"78",x"c0",x"48"),
    39 => (x"c0",x"4b",x"a6",x"e4"),
    40 => (x"48",x"49",x"66",x"e0"),
    41 => (x"e4",x"c0",x"80",x"c1"),
    42 => (x"48",x"11",x"58",x"a6"),
    43 => (x"70",x"58",x"a6",x"c4"),
    44 => (x"f6",x"c3",x"02",x"98"),
    45 => (x"02",x"66",x"c4",x"87"),
    46 => (x"c4",x"87",x"c6",x"c3"),
    47 => (x"78",x"c0",x"48",x"a6"),
    48 => (x"f0",x"c0",x"4a",x"6e"),
    49 => (x"da",x"c2",x"02",x"8a"),
    50 => (x"8a",x"f3",x"c0",x"87"),
    51 => (x"87",x"db",x"c2",x"02"),
    52 => (x"dc",x"02",x"8a",x"c1"),
    53 => (x"02",x"8a",x"c8",x"87"),
    54 => (x"c4",x"87",x"c8",x"c2"),
    55 => (x"87",x"d1",x"02",x"8a"),
    56 => (x"c1",x"02",x"8a",x"c3"),
    57 => (x"8a",x"c2",x"87",x"eb"),
    58 => (x"c3",x"87",x"c6",x"02"),
    59 => (x"c9",x"c2",x"05",x"8a"),
    60 => (x"73",x"83",x"c4",x"87"),
    61 => (x"69",x"89",x"c4",x"49"),
    62 => (x"c1",x"02",x"6e",x"7e"),
    63 => (x"a6",x"c8",x"87",x"c8"),
    64 => (x"c4",x"78",x"c0",x"48"),
    65 => (x"cc",x"78",x"c0",x"80"),
    66 => (x"4a",x"6e",x"4d",x"66"),
    67 => (x"cf",x"2a",x"b7",x"dc"),
    68 => (x"c4",x"48",x"6e",x"9a"),
    69 => (x"72",x"58",x"a6",x"30"),
    70 => (x"87",x"c5",x"02",x"9a"),
    71 => (x"c1",x"48",x"a6",x"c8"),
    72 => (x"06",x"aa",x"c9",x"78"),
    73 => (x"f7",x"c0",x"87",x"c5"),
    74 => (x"c0",x"87",x"c3",x"82"),
    75 => (x"66",x"c8",x"82",x"f0"),
    76 => (x"72",x"87",x"c7",x"02"),
    77 => (x"87",x"ff",x"c1",x"49"),
    78 => (x"85",x"c1",x"84",x"c1"),
    79 => (x"04",x"ad",x"b7",x"c8"),
    80 => (x"c1",x"87",x"c7",x"ff"),
    81 => (x"f0",x"c0",x"87",x"cf"),
    82 => (x"87",x"eb",x"c1",x"49"),
    83 => (x"c4",x"c1",x"84",x"c1"),
    84 => (x"73",x"83",x"c4",x"87"),
    85 => (x"6a",x"8a",x"c4",x"4a"),
    86 => (x"87",x"f7",x"c1",x"49"),
    87 => (x"4c",x"a4",x"49",x"70"),
    88 => (x"c4",x"87",x"f2",x"c0"),
    89 => (x"78",x"c1",x"48",x"a6"),
    90 => (x"c4",x"87",x"ea",x"c0"),
    91 => (x"c4",x"4a",x"73",x"83"),
    92 => (x"c1",x"49",x"6a",x"8a"),
    93 => (x"84",x"c1",x"87",x"c1"),
    94 => (x"49",x"6e",x"87",x"db"),
    95 => (x"d4",x"87",x"f8",x"c0"),
    96 => (x"c0",x"48",x"6e",x"87"),
    97 => (x"c7",x"05",x"a8",x"e5"),
    98 => (x"48",x"a6",x"c4",x"87"),
    99 => (x"87",x"c5",x"78",x"c1"),
   100 => (x"e2",x"c0",x"49",x"6e"),
   101 => (x"66",x"e0",x"c0",x"87"),
   102 => (x"80",x"c1",x"48",x"49"),
   103 => (x"58",x"a6",x"e4",x"c0"),
   104 => (x"a6",x"c4",x"48",x"11"),
   105 => (x"05",x"98",x"70",x"58"),
   106 => (x"74",x"87",x"ca",x"fc"),
   107 => (x"26",x"8e",x"f0",x"48"),
   108 => (x"26",x"4c",x"26",x"4d"),
   109 => (x"1e",x"4f",x"26",x"4b"),
   110 => (x"4a",x"71",x"86",x"fc"),
   111 => (x"69",x"49",x"c0",x"ff"),
   112 => (x"98",x"c0",x"c4",x"48"),
   113 => (x"70",x"58",x"a6",x"c4"),
   114 => (x"87",x"f3",x"02",x"98"),
   115 => (x"fc",x"48",x"79",x"72"),
   116 => (x"0e",x"4f",x"26",x"8e"),
   117 => (x"0e",x"5c",x"5b",x"5e"),
   118 => (x"4c",x"c0",x"4b",x"71"),
   119 => (x"02",x"9a",x"4a",x"13"),
   120 => (x"49",x"72",x"87",x"cd"),
   121 => (x"c1",x"87",x"d0",x"ff"),
   122 => (x"9a",x"4a",x"13",x"84"),
   123 => (x"74",x"87",x"f3",x"05"),
   124 => (x"26",x"4c",x"26",x"48"),
   125 => (x"1e",x"4f",x"26",x"4b"),
   126 => (x"1e",x"73",x"1e",x"72"),
   127 => (x"02",x"11",x"48",x"12"),
   128 => (x"c3",x"4b",x"87",x"ca"),
   129 => (x"73",x"9b",x"98",x"df"),
   130 => (x"87",x"f0",x"02",x"88"),
   131 => (x"4a",x"26",x"4b",x"26"),
   132 => (x"73",x"1e",x"4f",x"26"),
   133 => (x"c1",x"1e",x"72",x"1e"),
   134 => (x"87",x"ca",x"04",x"8b"),
   135 => (x"02",x"11",x"48",x"12"),
   136 => (x"02",x"88",x"87",x"c4"),
   137 => (x"4a",x"26",x"87",x"f1"),
   138 => (x"4f",x"26",x"4b",x"26"),
   139 => (x"81",x"48",x"73",x"1e"),
   140 => (x"c5",x"02",x"a9",x"73"),
   141 => (x"05",x"53",x"12",x"87"),
   142 => (x"4f",x"26",x"87",x"f6"),
   143 => (x"71",x"1e",x"73",x"1e"),
   144 => (x"4b",x"66",x"c8",x"4a"),
   145 => (x"71",x"8b",x"c1",x"49"),
   146 => (x"87",x"cf",x"02",x"99"),
   147 => (x"d4",x"ff",x"48",x"12"),
   148 => (x"49",x"73",x"78",x"08"),
   149 => (x"99",x"71",x"8b",x"c1"),
   150 => (x"26",x"87",x"f1",x"05"),
   151 => (x"0e",x"4f",x"26",x"4b"),
   152 => (x"0e",x"5c",x"5b",x"5e"),
   153 => (x"d4",x"ff",x"4a",x"71"),
   154 => (x"4b",x"66",x"cc",x"4c"),
   155 => (x"71",x"8b",x"c1",x"49"),
   156 => (x"87",x"ce",x"02",x"99"),
   157 => (x"6c",x"7c",x"ff",x"c3"),
   158 => (x"c1",x"49",x"73",x"52"),
   159 => (x"05",x"99",x"71",x"8b"),
   160 => (x"4c",x"26",x"87",x"f2"),
   161 => (x"4f",x"26",x"4b",x"26"),
   162 => (x"ff",x"1e",x"73",x"1e"),
   163 => (x"ff",x"c3",x"4b",x"d4"),
   164 => (x"c3",x"4a",x"6b",x"7b"),
   165 => (x"49",x"6b",x"7b",x"ff"),
   166 => (x"b1",x"72",x"32",x"c8"),
   167 => (x"6b",x"7b",x"ff",x"c3"),
   168 => (x"71",x"31",x"c8",x"4a"),
   169 => (x"7b",x"ff",x"c3",x"b2"),
   170 => (x"32",x"c8",x"49",x"6b"),
   171 => (x"48",x"71",x"b1",x"72"),
   172 => (x"4f",x"26",x"4b",x"26"),
   173 => (x"5c",x"5b",x"5e",x"0e"),
   174 => (x"4d",x"71",x"0e",x"5d"),
   175 => (x"75",x"4c",x"d4",x"ff"),
   176 => (x"98",x"ff",x"c3",x"48"),
   177 => (x"e8",x"c2",x"7c",x"70"),
   178 => (x"c8",x"05",x"bf",x"c0"),
   179 => (x"48",x"66",x"d0",x"87"),
   180 => (x"a6",x"d4",x"30",x"c9"),
   181 => (x"49",x"66",x"d0",x"58"),
   182 => (x"48",x"71",x"29",x"d8"),
   183 => (x"70",x"98",x"ff",x"c3"),
   184 => (x"49",x"66",x"d0",x"7c"),
   185 => (x"48",x"71",x"29",x"d0"),
   186 => (x"70",x"98",x"ff",x"c3"),
   187 => (x"49",x"66",x"d0",x"7c"),
   188 => (x"48",x"71",x"29",x"c8"),
   189 => (x"70",x"98",x"ff",x"c3"),
   190 => (x"48",x"66",x"d0",x"7c"),
   191 => (x"70",x"98",x"ff",x"c3"),
   192 => (x"d0",x"49",x"75",x"7c"),
   193 => (x"c3",x"48",x"71",x"29"),
   194 => (x"7c",x"70",x"98",x"ff"),
   195 => (x"f0",x"c9",x"4b",x"6c"),
   196 => (x"ff",x"c3",x"4a",x"ff"),
   197 => (x"87",x"cf",x"05",x"ab"),
   198 => (x"6c",x"7c",x"71",x"49"),
   199 => (x"02",x"8a",x"c1",x"4b"),
   200 => (x"ab",x"71",x"87",x"c5"),
   201 => (x"73",x"87",x"f2",x"02"),
   202 => (x"26",x"4d",x"26",x"48"),
   203 => (x"26",x"4b",x"26",x"4c"),
   204 => (x"49",x"c0",x"1e",x"4f"),
   205 => (x"c3",x"48",x"d4",x"ff"),
   206 => (x"81",x"c1",x"78",x"ff"),
   207 => (x"a9",x"b7",x"c8",x"c3"),
   208 => (x"26",x"87",x"f1",x"04"),
   209 => (x"5b",x"5e",x"0e",x"4f"),
   210 => (x"c0",x"0e",x"5d",x"5c"),
   211 => (x"f7",x"c1",x"f0",x"ff"),
   212 => (x"c0",x"c0",x"c1",x"4d"),
   213 => (x"4b",x"c0",x"c0",x"c0"),
   214 => (x"c4",x"87",x"d6",x"ff"),
   215 => (x"c0",x"4c",x"df",x"f8"),
   216 => (x"fd",x"49",x"75",x"1e"),
   217 => (x"86",x"c4",x"87",x"ce"),
   218 => (x"c0",x"05",x"a8",x"c1"),
   219 => (x"d4",x"ff",x"87",x"e5"),
   220 => (x"78",x"ff",x"c3",x"48"),
   221 => (x"e1",x"c0",x"1e",x"73"),
   222 => (x"49",x"e9",x"c1",x"f0"),
   223 => (x"c4",x"87",x"f5",x"fc"),
   224 => (x"05",x"98",x"70",x"86"),
   225 => (x"d4",x"ff",x"87",x"ca"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"87",x"cb",x"48",x"c1"),
   228 => (x"c1",x"87",x"de",x"fe"),
   229 => (x"c6",x"ff",x"05",x"8c"),
   230 => (x"26",x"48",x"c0",x"87"),
   231 => (x"26",x"4c",x"26",x"4d"),
   232 => (x"0e",x"4f",x"26",x"4b"),
   233 => (x"0e",x"5c",x"5b",x"5e"),
   234 => (x"c1",x"f0",x"ff",x"c0"),
   235 => (x"d4",x"ff",x"4c",x"c1"),
   236 => (x"78",x"ff",x"c3",x"48"),
   237 => (x"f8",x"49",x"e8",x"cf"),
   238 => (x"4b",x"d3",x"87",x"d9"),
   239 => (x"49",x"74",x"1e",x"c0"),
   240 => (x"c4",x"87",x"f1",x"fb"),
   241 => (x"05",x"98",x"70",x"86"),
   242 => (x"d4",x"ff",x"87",x"ca"),
   243 => (x"78",x"ff",x"c3",x"48"),
   244 => (x"87",x"cb",x"48",x"c1"),
   245 => (x"c1",x"87",x"da",x"fd"),
   246 => (x"df",x"ff",x"05",x"8b"),
   247 => (x"26",x"48",x"c0",x"87"),
   248 => (x"26",x"4b",x"26",x"4c"),
   249 => (x"00",x"00",x"00",x"4f"),
   250 => (x"00",x"44",x"4d",x"43"),
   251 => (x"43",x"48",x"44",x"53"),
   252 => (x"69",x"61",x"66",x"20"),
   253 => (x"00",x"0a",x"21",x"6c"),
   254 => (x"52",x"52",x"45",x"49"),
   255 => (x"00",x"00",x"00",x"00"),
   256 => (x"00",x"49",x"50",x"53"),
   257 => (x"74",x"69",x"72",x"57"),
   258 => (x"61",x"66",x"20",x"65"),
   259 => (x"64",x"65",x"6c",x"69"),
   260 => (x"5e",x"0e",x"00",x"0a"),
   261 => (x"0e",x"5d",x"5c",x"5b"),
   262 => (x"ff",x"4d",x"ff",x"c3"),
   263 => (x"d0",x"fc",x"4b",x"d4"),
   264 => (x"1e",x"ea",x"c6",x"87"),
   265 => (x"c1",x"f0",x"e1",x"c0"),
   266 => (x"c7",x"fa",x"49",x"c8"),
   267 => (x"c1",x"86",x"c4",x"87"),
   268 => (x"87",x"c8",x"02",x"a8"),
   269 => (x"c0",x"87",x"ec",x"fd"),
   270 => (x"87",x"e8",x"c1",x"48"),
   271 => (x"70",x"87",x"c9",x"f9"),
   272 => (x"ff",x"ff",x"cf",x"49"),
   273 => (x"a9",x"ea",x"c6",x"99"),
   274 => (x"fd",x"87",x"c8",x"02"),
   275 => (x"48",x"c0",x"87",x"d5"),
   276 => (x"75",x"87",x"d1",x"c1"),
   277 => (x"4c",x"f1",x"c0",x"7b"),
   278 => (x"70",x"87",x"ea",x"fb"),
   279 => (x"ec",x"c0",x"02",x"98"),
   280 => (x"c0",x"1e",x"c0",x"87"),
   281 => (x"fa",x"c1",x"f0",x"ff"),
   282 => (x"87",x"c8",x"f9",x"49"),
   283 => (x"98",x"70",x"86",x"c4"),
   284 => (x"75",x"87",x"da",x"05"),
   285 => (x"75",x"49",x"6b",x"7b"),
   286 => (x"75",x"7b",x"75",x"7b"),
   287 => (x"c1",x"7b",x"75",x"7b"),
   288 => (x"c4",x"02",x"99",x"c0"),
   289 => (x"db",x"48",x"c1",x"87"),
   290 => (x"d7",x"48",x"c0",x"87"),
   291 => (x"05",x"ac",x"c2",x"87"),
   292 => (x"ec",x"cf",x"87",x"ca"),
   293 => (x"87",x"fb",x"f4",x"49"),
   294 => (x"87",x"c8",x"48",x"c0"),
   295 => (x"fe",x"05",x"8c",x"c1"),
   296 => (x"48",x"c0",x"87",x"f6"),
   297 => (x"4c",x"26",x"4d",x"26"),
   298 => (x"4f",x"26",x"4b",x"26"),
   299 => (x"5c",x"5b",x"5e",x"0e"),
   300 => (x"d0",x"ff",x"0e",x"5d"),
   301 => (x"d0",x"e5",x"c0",x"4d"),
   302 => (x"c2",x"4c",x"c0",x"c1"),
   303 => (x"c1",x"48",x"c0",x"e8"),
   304 => (x"49",x"c0",x"d0",x"78"),
   305 => (x"c7",x"87",x"cc",x"f4"),
   306 => (x"f9",x"7d",x"c2",x"4b"),
   307 => (x"7d",x"c3",x"87",x"e3"),
   308 => (x"49",x"74",x"1e",x"c0"),
   309 => (x"c4",x"87",x"dd",x"f7"),
   310 => (x"05",x"a8",x"c1",x"86"),
   311 => (x"c2",x"4b",x"87",x"c1"),
   312 => (x"87",x"cb",x"05",x"ab"),
   313 => (x"f3",x"49",x"f8",x"cf"),
   314 => (x"48",x"c0",x"87",x"e9"),
   315 => (x"c1",x"87",x"f6",x"c0"),
   316 => (x"d4",x"ff",x"05",x"8b"),
   317 => (x"87",x"da",x"fc",x"87"),
   318 => (x"58",x"c4",x"e8",x"c2"),
   319 => (x"cd",x"05",x"98",x"70"),
   320 => (x"c0",x"1e",x"c1",x"87"),
   321 => (x"d0",x"c1",x"f0",x"ff"),
   322 => (x"87",x"e8",x"f6",x"49"),
   323 => (x"d4",x"ff",x"86",x"c4"),
   324 => (x"78",x"ff",x"c3",x"48"),
   325 => (x"c2",x"87",x"ee",x"c4"),
   326 => (x"c2",x"58",x"c8",x"e8"),
   327 => (x"48",x"d4",x"ff",x"7d"),
   328 => (x"c1",x"78",x"ff",x"c3"),
   329 => (x"26",x"4d",x"26",x"48"),
   330 => (x"26",x"4b",x"26",x"4c"),
   331 => (x"5b",x"5e",x"0e",x"4f"),
   332 => (x"71",x"0e",x"5d",x"5c"),
   333 => (x"4c",x"ff",x"c3",x"4d"),
   334 => (x"74",x"4b",x"d4",x"ff"),
   335 => (x"48",x"d0",x"ff",x"7b"),
   336 => (x"74",x"78",x"c3",x"c4"),
   337 => (x"c0",x"1e",x"75",x"7b"),
   338 => (x"d8",x"c1",x"f0",x"ff"),
   339 => (x"87",x"e4",x"f5",x"49"),
   340 => (x"98",x"70",x"86",x"c4"),
   341 => (x"d0",x"87",x"cb",x"02"),
   342 => (x"f6",x"f1",x"49",x"c4"),
   343 => (x"c0",x"48",x"c1",x"87"),
   344 => (x"7b",x"74",x"87",x"ee"),
   345 => (x"c8",x"7b",x"fe",x"c3"),
   346 => (x"66",x"d4",x"1e",x"c0"),
   347 => (x"87",x"cc",x"f3",x"49"),
   348 => (x"7b",x"74",x"86",x"c4"),
   349 => (x"7b",x"74",x"7b",x"74"),
   350 => (x"4a",x"e0",x"da",x"d8"),
   351 => (x"05",x"6b",x"7b",x"74"),
   352 => (x"8a",x"c1",x"87",x"c5"),
   353 => (x"74",x"87",x"f5",x"05"),
   354 => (x"48",x"d0",x"ff",x"7b"),
   355 => (x"48",x"c0",x"78",x"c2"),
   356 => (x"4c",x"26",x"4d",x"26"),
   357 => (x"4f",x"26",x"4b",x"26"),
   358 => (x"5c",x"5b",x"5e",x"0e"),
   359 => (x"86",x"fc",x"0e",x"5d"),
   360 => (x"d4",x"ff",x"4b",x"71"),
   361 => (x"c5",x"7e",x"c0",x"4c"),
   362 => (x"4a",x"df",x"cd",x"ee"),
   363 => (x"6c",x"7c",x"ff",x"c3"),
   364 => (x"a8",x"fe",x"c3",x"48"),
   365 => (x"87",x"f8",x"c0",x"05"),
   366 => (x"9b",x"73",x"4d",x"74"),
   367 => (x"d4",x"87",x"cc",x"02"),
   368 => (x"49",x"73",x"1e",x"66"),
   369 => (x"c4",x"87",x"d8",x"f2"),
   370 => (x"ff",x"87",x"d4",x"86"),
   371 => (x"d1",x"c4",x"48",x"d0"),
   372 => (x"4a",x"66",x"d4",x"78"),
   373 => (x"c1",x"7d",x"ff",x"c3"),
   374 => (x"87",x"f8",x"05",x"8a"),
   375 => (x"c3",x"5a",x"a6",x"d8"),
   376 => (x"73",x"7c",x"7c",x"ff"),
   377 => (x"87",x"c5",x"05",x"9b"),
   378 => (x"d0",x"48",x"d0",x"ff"),
   379 => (x"7e",x"4a",x"c1",x"78"),
   380 => (x"fe",x"05",x"8a",x"c1"),
   381 => (x"48",x"6e",x"87",x"f6"),
   382 => (x"4d",x"26",x"8e",x"fc"),
   383 => (x"4b",x"26",x"4c",x"26"),
   384 => (x"73",x"1e",x"4f",x"26"),
   385 => (x"c0",x"4a",x"71",x"1e"),
   386 => (x"48",x"d4",x"ff",x"4b"),
   387 => (x"ff",x"78",x"ff",x"c3"),
   388 => (x"c3",x"c4",x"48",x"d0"),
   389 => (x"48",x"d4",x"ff",x"78"),
   390 => (x"72",x"78",x"ff",x"c3"),
   391 => (x"f0",x"ff",x"c0",x"1e"),
   392 => (x"f2",x"49",x"d1",x"c1"),
   393 => (x"86",x"c4",x"87",x"ce"),
   394 => (x"d2",x"05",x"98",x"70"),
   395 => (x"1e",x"c0",x"c8",x"87"),
   396 => (x"fd",x"49",x"66",x"cc"),
   397 => (x"86",x"c4",x"87",x"e2"),
   398 => (x"d0",x"ff",x"4b",x"70"),
   399 => (x"73",x"78",x"c2",x"48"),
   400 => (x"26",x"4b",x"26",x"48"),
   401 => (x"5b",x"5e",x"0e",x"4f"),
   402 => (x"c0",x"0e",x"5d",x"5c"),
   403 => (x"f0",x"ff",x"c0",x"1e"),
   404 => (x"f1",x"49",x"c9",x"c1"),
   405 => (x"1e",x"d2",x"87",x"de"),
   406 => (x"49",x"d0",x"e8",x"c2"),
   407 => (x"c8",x"87",x"f9",x"fc"),
   408 => (x"c1",x"4c",x"c0",x"86"),
   409 => (x"ac",x"b7",x"d2",x"84"),
   410 => (x"c2",x"87",x"f8",x"04"),
   411 => (x"bf",x"97",x"d0",x"e8"),
   412 => (x"99",x"c0",x"c3",x"49"),
   413 => (x"05",x"a9",x"c0",x"c1"),
   414 => (x"c2",x"87",x"e7",x"c0"),
   415 => (x"bf",x"97",x"d7",x"e8"),
   416 => (x"c2",x"31",x"d0",x"49"),
   417 => (x"bf",x"97",x"d8",x"e8"),
   418 => (x"72",x"32",x"c8",x"4a"),
   419 => (x"d9",x"e8",x"c2",x"b1"),
   420 => (x"b1",x"4a",x"bf",x"97"),
   421 => (x"ff",x"cf",x"4c",x"71"),
   422 => (x"c1",x"9c",x"ff",x"ff"),
   423 => (x"c1",x"34",x"ca",x"84"),
   424 => (x"e8",x"c2",x"87",x"e7"),
   425 => (x"49",x"bf",x"97",x"d9"),
   426 => (x"99",x"c6",x"31",x"c1"),
   427 => (x"97",x"da",x"e8",x"c2"),
   428 => (x"b7",x"c7",x"4a",x"bf"),
   429 => (x"c2",x"b1",x"72",x"2a"),
   430 => (x"bf",x"97",x"d5",x"e8"),
   431 => (x"9d",x"cf",x"4d",x"4a"),
   432 => (x"97",x"d6",x"e8",x"c2"),
   433 => (x"9a",x"c3",x"4a",x"bf"),
   434 => (x"e8",x"c2",x"32",x"ca"),
   435 => (x"4b",x"bf",x"97",x"d7"),
   436 => (x"b2",x"73",x"33",x"c2"),
   437 => (x"97",x"d8",x"e8",x"c2"),
   438 => (x"c0",x"c3",x"4b",x"bf"),
   439 => (x"2b",x"b7",x"c6",x"9b"),
   440 => (x"81",x"c2",x"b2",x"73"),
   441 => (x"30",x"71",x"48",x"c1"),
   442 => (x"48",x"c1",x"49",x"70"),
   443 => (x"4d",x"70",x"30",x"75"),
   444 => (x"84",x"c1",x"4c",x"72"),
   445 => (x"c0",x"c8",x"94",x"71"),
   446 => (x"cc",x"06",x"ad",x"b7"),
   447 => (x"b7",x"34",x"c1",x"87"),
   448 => (x"b7",x"c0",x"c8",x"2d"),
   449 => (x"f4",x"ff",x"01",x"ad"),
   450 => (x"26",x"48",x"74",x"87"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"0e",x"4f",x"26",x"4b"),
   453 => (x"5d",x"5c",x"5b",x"5e"),
   454 => (x"c2",x"86",x"fc",x"0e"),
   455 => (x"c0",x"48",x"f8",x"f0"),
   456 => (x"f0",x"e8",x"c2",x"78"),
   457 => (x"fb",x"49",x"c0",x"1e"),
   458 => (x"86",x"c4",x"87",x"d8"),
   459 => (x"c5",x"05",x"98",x"70"),
   460 => (x"c9",x"48",x"c0",x"87"),
   461 => (x"4d",x"c0",x"87",x"d7"),
   462 => (x"48",x"f4",x"f5",x"c2"),
   463 => (x"e9",x"c2",x"78",x"c1"),
   464 => (x"e6",x"c0",x"4a",x"e6"),
   465 => (x"4b",x"c8",x"49",x"e4"),
   466 => (x"70",x"87",x"c7",x"eb"),
   467 => (x"87",x"c6",x"05",x"98"),
   468 => (x"48",x"f4",x"f5",x"c2"),
   469 => (x"ea",x"c2",x"78",x"c0"),
   470 => (x"e6",x"c0",x"4a",x"c2"),
   471 => (x"4b",x"c8",x"49",x"f0"),
   472 => (x"70",x"87",x"ef",x"ea"),
   473 => (x"87",x"c6",x"05",x"98"),
   474 => (x"48",x"f4",x"f5",x"c2"),
   475 => (x"f5",x"c2",x"78",x"c0"),
   476 => (x"c0",x"02",x"bf",x"f4"),
   477 => (x"ef",x"c2",x"87",x"ff"),
   478 => (x"c2",x"4d",x"bf",x"f6"),
   479 => (x"bf",x"9f",x"ee",x"f0"),
   480 => (x"58",x"a6",x"c4",x"48"),
   481 => (x"a8",x"ea",x"d6",x"c5"),
   482 => (x"c2",x"87",x"c7",x"05"),
   483 => (x"4d",x"bf",x"f6",x"ef"),
   484 => (x"48",x"6e",x"87",x"ce"),
   485 => (x"a8",x"d5",x"e9",x"ca"),
   486 => (x"c0",x"87",x"c5",x"02"),
   487 => (x"87",x"ed",x"c7",x"48"),
   488 => (x"1e",x"f0",x"e8",x"c2"),
   489 => (x"d9",x"f9",x"49",x"75"),
   490 => (x"70",x"86",x"c4",x"87"),
   491 => (x"87",x"c5",x"05",x"98"),
   492 => (x"d8",x"c7",x"48",x"c0"),
   493 => (x"c2",x"ea",x"c2",x"87"),
   494 => (x"fc",x"e6",x"c0",x"4a"),
   495 => (x"e9",x"4b",x"c8",x"49"),
   496 => (x"98",x"70",x"87",x"d0"),
   497 => (x"87",x"c8",x"c0",x"05"),
   498 => (x"48",x"f8",x"f0",x"c2"),
   499 => (x"87",x"d8",x"78",x"c1"),
   500 => (x"4a",x"e6",x"e9",x"c2"),
   501 => (x"49",x"c8",x"e7",x"c0"),
   502 => (x"f5",x"e8",x"4b",x"c8"),
   503 => (x"02",x"98",x"70",x"87"),
   504 => (x"c0",x"87",x"c5",x"c0"),
   505 => (x"87",x"e5",x"c6",x"48"),
   506 => (x"97",x"ee",x"f0",x"c2"),
   507 => (x"d5",x"c1",x"49",x"bf"),
   508 => (x"cd",x"c0",x"05",x"a9"),
   509 => (x"ef",x"f0",x"c2",x"87"),
   510 => (x"c2",x"49",x"bf",x"97"),
   511 => (x"c0",x"02",x"a9",x"ea"),
   512 => (x"48",x"c0",x"87",x"c5"),
   513 => (x"c2",x"87",x"c6",x"c6"),
   514 => (x"bf",x"97",x"f0",x"e8"),
   515 => (x"58",x"a6",x"c4",x"48"),
   516 => (x"02",x"a8",x"e9",x"c3"),
   517 => (x"6e",x"87",x"ce",x"c0"),
   518 => (x"a8",x"eb",x"c3",x"48"),
   519 => (x"87",x"c5",x"c0",x"02"),
   520 => (x"e8",x"c5",x"48",x"c0"),
   521 => (x"fb",x"e8",x"c2",x"87"),
   522 => (x"99",x"49",x"bf",x"97"),
   523 => (x"87",x"cc",x"c0",x"05"),
   524 => (x"97",x"fc",x"e8",x"c2"),
   525 => (x"a9",x"c2",x"49",x"bf"),
   526 => (x"87",x"c5",x"c0",x"02"),
   527 => (x"cc",x"c5",x"48",x"c0"),
   528 => (x"fd",x"e8",x"c2",x"87"),
   529 => (x"c2",x"48",x"bf",x"97"),
   530 => (x"70",x"58",x"f4",x"f0"),
   531 => (x"88",x"c1",x"48",x"4c"),
   532 => (x"58",x"f8",x"f0",x"c2"),
   533 => (x"97",x"fe",x"e8",x"c2"),
   534 => (x"81",x"75",x"49",x"bf"),
   535 => (x"97",x"ff",x"e8",x"c2"),
   536 => (x"32",x"c8",x"4a",x"bf"),
   537 => (x"c2",x"7e",x"a1",x"72"),
   538 => (x"6e",x"48",x"d0",x"f5"),
   539 => (x"c0",x"e9",x"c2",x"78"),
   540 => (x"c2",x"48",x"bf",x"97"),
   541 => (x"c2",x"58",x"e8",x"f5"),
   542 => (x"02",x"bf",x"f8",x"f0"),
   543 => (x"c2",x"87",x"d3",x"c2"),
   544 => (x"c0",x"4a",x"c2",x"ea"),
   545 => (x"c8",x"49",x"d8",x"e6"),
   546 => (x"87",x"c6",x"e6",x"4b"),
   547 => (x"c0",x"02",x"98",x"70"),
   548 => (x"48",x"c0",x"87",x"c5"),
   549 => (x"c2",x"87",x"f6",x"c3"),
   550 => (x"4c",x"bf",x"f0",x"f0"),
   551 => (x"5c",x"e4",x"f5",x"c2"),
   552 => (x"97",x"d5",x"e9",x"c2"),
   553 => (x"31",x"c8",x"49",x"bf"),
   554 => (x"97",x"d4",x"e9",x"c2"),
   555 => (x"49",x"a1",x"4a",x"bf"),
   556 => (x"97",x"d6",x"e9",x"c2"),
   557 => (x"32",x"d0",x"4a",x"bf"),
   558 => (x"c2",x"49",x"a1",x"72"),
   559 => (x"bf",x"97",x"d7",x"e9"),
   560 => (x"72",x"32",x"d8",x"4a"),
   561 => (x"f5",x"c2",x"49",x"a1"),
   562 => (x"f5",x"c2",x"59",x"ec"),
   563 => (x"c2",x"91",x"bf",x"e4"),
   564 => (x"81",x"bf",x"d0",x"f5"),
   565 => (x"59",x"d8",x"f5",x"c2"),
   566 => (x"97",x"dd",x"e9",x"c2"),
   567 => (x"32",x"c8",x"4a",x"bf"),
   568 => (x"97",x"dc",x"e9",x"c2"),
   569 => (x"4a",x"a2",x"4b",x"bf"),
   570 => (x"97",x"de",x"e9",x"c2"),
   571 => (x"33",x"d0",x"4b",x"bf"),
   572 => (x"c2",x"4a",x"a2",x"73"),
   573 => (x"bf",x"97",x"df",x"e9"),
   574 => (x"d8",x"9b",x"cf",x"4b"),
   575 => (x"4a",x"a2",x"73",x"33"),
   576 => (x"5a",x"dc",x"f5",x"c2"),
   577 => (x"92",x"74",x"8a",x"c2"),
   578 => (x"48",x"dc",x"f5",x"c2"),
   579 => (x"c1",x"78",x"a1",x"72"),
   580 => (x"e9",x"c2",x"87",x"c7"),
   581 => (x"49",x"bf",x"97",x"c2"),
   582 => (x"e9",x"c2",x"31",x"c8"),
   583 => (x"4a",x"bf",x"97",x"c1"),
   584 => (x"31",x"c5",x"49",x"a1"),
   585 => (x"c9",x"81",x"ff",x"c7"),
   586 => (x"e4",x"f5",x"c2",x"29"),
   587 => (x"c7",x"e9",x"c2",x"59"),
   588 => (x"c8",x"4a",x"bf",x"97"),
   589 => (x"c6",x"e9",x"c2",x"32"),
   590 => (x"a2",x"4b",x"bf",x"97"),
   591 => (x"ec",x"f5",x"c2",x"4a"),
   592 => (x"e4",x"f5",x"c2",x"5a"),
   593 => (x"82",x"6e",x"92",x"bf"),
   594 => (x"5a",x"e0",x"f5",x"c2"),
   595 => (x"48",x"d8",x"f5",x"c2"),
   596 => (x"f5",x"c2",x"78",x"c0"),
   597 => (x"a1",x"72",x"48",x"d4"),
   598 => (x"ec",x"f5",x"c2",x"78"),
   599 => (x"d8",x"f5",x"c2",x"48"),
   600 => (x"f5",x"c2",x"78",x"bf"),
   601 => (x"f5",x"c2",x"48",x"f0"),
   602 => (x"c2",x"78",x"bf",x"dc"),
   603 => (x"02",x"bf",x"f8",x"f0"),
   604 => (x"74",x"87",x"c9",x"c0"),
   605 => (x"a6",x"30",x"c4",x"48"),
   606 => (x"87",x"c9",x"c0",x"58"),
   607 => (x"bf",x"e0",x"f5",x"c2"),
   608 => (x"a6",x"30",x"c4",x"48"),
   609 => (x"fc",x"f0",x"c2",x"58"),
   610 => (x"c1",x"78",x"6e",x"48"),
   611 => (x"26",x"8e",x"fc",x"48"),
   612 => (x"26",x"4c",x"26",x"4d"),
   613 => (x"00",x"4f",x"26",x"4b"),
   614 => (x"33",x"54",x"41",x"46"),
   615 => (x"20",x"20",x"20",x"32"),
   616 => (x"00",x"00",x"00",x"00"),
   617 => (x"31",x"54",x"41",x"46"),
   618 => (x"20",x"20",x"20",x"36"),
   619 => (x"00",x"00",x"00",x"00"),
   620 => (x"33",x"54",x"41",x"46"),
   621 => (x"20",x"20",x"20",x"32"),
   622 => (x"00",x"00",x"00",x"00"),
   623 => (x"33",x"54",x"41",x"46"),
   624 => (x"20",x"20",x"20",x"32"),
   625 => (x"00",x"00",x"00",x"00"),
   626 => (x"31",x"54",x"41",x"46"),
   627 => (x"20",x"20",x"20",x"36"),
   628 => (x"5b",x"5e",x"0e",x"00"),
   629 => (x"71",x"0e",x"5d",x"5c"),
   630 => (x"f8",x"f0",x"c2",x"4a"),
   631 => (x"87",x"cb",x"02",x"bf"),
   632 => (x"2b",x"c7",x"4b",x"72"),
   633 => (x"ff",x"c1",x"4d",x"72"),
   634 => (x"72",x"87",x"c9",x"9d"),
   635 => (x"72",x"2b",x"c8",x"4b"),
   636 => (x"9d",x"ff",x"c3",x"4d"),
   637 => (x"bf",x"d0",x"f5",x"c2"),
   638 => (x"dc",x"fe",x"c0",x"83"),
   639 => (x"d9",x"02",x"ab",x"bf"),
   640 => (x"e0",x"fe",x"c0",x"87"),
   641 => (x"f0",x"e8",x"c2",x"5b"),
   642 => (x"ef",x"49",x"73",x"1e"),
   643 => (x"86",x"c4",x"87",x"f4"),
   644 => (x"c5",x"05",x"98",x"70"),
   645 => (x"c0",x"48",x"c0",x"87"),
   646 => (x"f0",x"c2",x"87",x"e6"),
   647 => (x"d2",x"02",x"bf",x"f8"),
   648 => (x"c4",x"49",x"75",x"87"),
   649 => (x"f0",x"e8",x"c2",x"91"),
   650 => (x"cf",x"4c",x"69",x"81"),
   651 => (x"ff",x"ff",x"ff",x"ff"),
   652 => (x"75",x"87",x"cb",x"9c"),
   653 => (x"c2",x"91",x"c2",x"49"),
   654 => (x"9f",x"81",x"f0",x"e8"),
   655 => (x"48",x"74",x"4c",x"69"),
   656 => (x"4c",x"26",x"4d",x"26"),
   657 => (x"4f",x"26",x"4b",x"26"),
   658 => (x"5c",x"5b",x"5e",x"0e"),
   659 => (x"86",x"f4",x"0e",x"5d"),
   660 => (x"c4",x"59",x"a6",x"c8"),
   661 => (x"80",x"c8",x"48",x"66"),
   662 => (x"6e",x"58",x"a6",x"c4"),
   663 => (x"1e",x"78",x"c0",x"48"),
   664 => (x"ff",x"cc",x"49",x"c1"),
   665 => (x"70",x"86",x"c4",x"87"),
   666 => (x"c0",x"02",x"9c",x"4c"),
   667 => (x"f1",x"c2",x"87",x"fc"),
   668 => (x"66",x"dc",x"4a",x"c0"),
   669 => (x"fe",x"dd",x"ff",x"49"),
   670 => (x"02",x"98",x"70",x"87"),
   671 => (x"74",x"87",x"eb",x"c0"),
   672 => (x"49",x"66",x"dc",x"4a"),
   673 => (x"de",x"ff",x"4b",x"cb"),
   674 => (x"98",x"70",x"87",x"c8"),
   675 => (x"c0",x"87",x"db",x"02"),
   676 => (x"02",x"9c",x"74",x"1e"),
   677 => (x"4d",x"c0",x"87",x"c4"),
   678 => (x"4d",x"c1",x"87",x"c2"),
   679 => (x"c3",x"cc",x"49",x"75"),
   680 => (x"70",x"86",x"c4",x"87"),
   681 => (x"ff",x"05",x"9c",x"4c"),
   682 => (x"9c",x"74",x"87",x"c4"),
   683 => (x"87",x"f5",x"c1",x"02"),
   684 => (x"6e",x"49",x"a4",x"dc"),
   685 => (x"da",x"78",x"69",x"48"),
   686 => (x"66",x"c4",x"49",x"a4"),
   687 => (x"9f",x"85",x"c4",x"4d"),
   688 => (x"f0",x"c2",x"7d",x"69"),
   689 => (x"d3",x"02",x"bf",x"f8"),
   690 => (x"49",x"a4",x"d4",x"87"),
   691 => (x"c0",x"49",x"69",x"9f"),
   692 => (x"71",x"99",x"ff",x"ff"),
   693 => (x"c4",x"30",x"d0",x"48"),
   694 => (x"87",x"c2",x"58",x"a6"),
   695 => (x"49",x"6e",x"7e",x"c0"),
   696 => (x"70",x"80",x"6d",x"48"),
   697 => (x"48",x"66",x"c4",x"7d"),
   698 => (x"66",x"c4",x"78",x"c0"),
   699 => (x"6d",x"81",x"cc",x"49"),
   700 => (x"49",x"66",x"c4",x"79"),
   701 => (x"79",x"c0",x"81",x"d0"),
   702 => (x"c0",x"48",x"a6",x"c8"),
   703 => (x"4c",x"66",x"c8",x"78"),
   704 => (x"d4",x"4a",x"66",x"c4"),
   705 => (x"c8",x"49",x"74",x"82"),
   706 => (x"49",x"a1",x"72",x"91"),
   707 => (x"79",x"6d",x"41",x"c0"),
   708 => (x"b7",x"c6",x"84",x"c1"),
   709 => (x"e7",x"ff",x"04",x"ac"),
   710 => (x"49",x"66",x"c4",x"87"),
   711 => (x"c0",x"81",x"c4",x"c1"),
   712 => (x"c2",x"48",x"c1",x"79"),
   713 => (x"f4",x"48",x"c0",x"87"),
   714 => (x"26",x"4d",x"26",x"8e"),
   715 => (x"26",x"4b",x"26",x"4c"),
   716 => (x"5b",x"5e",x"0e",x"4f"),
   717 => (x"71",x"0e",x"5d",x"5c"),
   718 => (x"4d",x"66",x"d0",x"4c"),
   719 => (x"75",x"85",x"49",x"6c"),
   720 => (x"f4",x"f0",x"c2",x"b9"),
   721 => (x"ba",x"ff",x"4a",x"bf"),
   722 => (x"99",x"71",x"99",x"72"),
   723 => (x"87",x"e4",x"c0",x"02"),
   724 => (x"6b",x"4b",x"a4",x"c4"),
   725 => (x"87",x"f9",x"f9",x"49"),
   726 => (x"f0",x"c2",x"7b",x"70"),
   727 => (x"6c",x"49",x"bf",x"f0"),
   728 => (x"75",x"7c",x"71",x"81"),
   729 => (x"f4",x"f0",x"c2",x"b9"),
   730 => (x"ba",x"ff",x"4a",x"bf"),
   731 => (x"99",x"71",x"99",x"72"),
   732 => (x"87",x"dc",x"ff",x"05"),
   733 => (x"4d",x"26",x"7c",x"75"),
   734 => (x"4b",x"26",x"4c",x"26"),
   735 => (x"73",x"1e",x"4f",x"26"),
   736 => (x"c2",x"4b",x"71",x"1e"),
   737 => (x"49",x"bf",x"d4",x"f5"),
   738 => (x"6a",x"4a",x"a3",x"c4"),
   739 => (x"c2",x"8a",x"c2",x"4a"),
   740 => (x"92",x"bf",x"f0",x"f0"),
   741 => (x"c2",x"49",x"a1",x"72"),
   742 => (x"4a",x"bf",x"f4",x"f0"),
   743 => (x"a1",x"72",x"9a",x"6b"),
   744 => (x"e0",x"fe",x"c0",x"49"),
   745 => (x"1e",x"66",x"c8",x"59"),
   746 => (x"87",x"d6",x"e9",x"71"),
   747 => (x"98",x"70",x"86",x"c4"),
   748 => (x"c0",x"87",x"c4",x"05"),
   749 => (x"c1",x"87",x"c2",x"48"),
   750 => (x"26",x"4b",x"26",x"48"),
   751 => (x"1e",x"73",x"1e",x"4f"),
   752 => (x"f5",x"c2",x"4b",x"71"),
   753 => (x"c4",x"49",x"bf",x"d4"),
   754 => (x"4a",x"6a",x"4a",x"a3"),
   755 => (x"f0",x"c2",x"8a",x"c2"),
   756 => (x"72",x"92",x"bf",x"f0"),
   757 => (x"f0",x"c2",x"49",x"a1"),
   758 => (x"6b",x"4a",x"bf",x"f4"),
   759 => (x"49",x"a1",x"72",x"9a"),
   760 => (x"59",x"e0",x"fe",x"c0"),
   761 => (x"71",x"1e",x"66",x"c8"),
   762 => (x"c4",x"87",x"c2",x"e5"),
   763 => (x"05",x"98",x"70",x"86"),
   764 => (x"48",x"c0",x"87",x"c4"),
   765 => (x"48",x"c1",x"87",x"c2"),
   766 => (x"4f",x"26",x"4b",x"26"),
   767 => (x"5c",x"5b",x"5e",x"0e"),
   768 => (x"86",x"e4",x"0e",x"5d"),
   769 => (x"ec",x"c0",x"4b",x"71"),
   770 => (x"28",x"c9",x"48",x"66"),
   771 => (x"c2",x"58",x"a6",x"cc"),
   772 => (x"49",x"bf",x"f4",x"f0"),
   773 => (x"48",x"71",x"b9",x"ff"),
   774 => (x"d4",x"98",x"66",x"c8"),
   775 => (x"48",x"71",x"58",x"a6"),
   776 => (x"a6",x"d0",x"98",x"6b"),
   777 => (x"7e",x"a3",x"c4",x"58"),
   778 => (x"6e",x"48",x"a6",x"c4"),
   779 => (x"66",x"d0",x"78",x"bf"),
   780 => (x"a8",x"66",x"cc",x"48"),
   781 => (x"c8",x"87",x"c6",x"05"),
   782 => (x"c7",x"c3",x"7b",x"66"),
   783 => (x"48",x"a6",x"d4",x"87"),
   784 => (x"ff",x"ff",x"ff",x"c1"),
   785 => (x"c4",x"78",x"ff",x"ff"),
   786 => (x"c0",x"78",x"ff",x"80"),
   787 => (x"4d",x"a3",x"d4",x"4a"),
   788 => (x"91",x"c8",x"49",x"72"),
   789 => (x"d0",x"49",x"a1",x"75"),
   790 => (x"8c",x"69",x"4c",x"66"),
   791 => (x"04",x"ac",x"b7",x"c0"),
   792 => (x"66",x"d4",x"87",x"cd"),
   793 => (x"c6",x"03",x"ac",x"b7"),
   794 => (x"5a",x"a6",x"dc",x"87"),
   795 => (x"c1",x"5c",x"a6",x"d8"),
   796 => (x"aa",x"b7",x"c6",x"82"),
   797 => (x"87",x"d5",x"ff",x"04"),
   798 => (x"c0",x"48",x"66",x"d8"),
   799 => (x"d0",x"04",x"a8",x"b7"),
   800 => (x"49",x"66",x"d8",x"87"),
   801 => (x"a1",x"75",x"91",x"c8"),
   802 => (x"6e",x"7b",x"21",x"49"),
   803 => (x"c9",x"78",x"69",x"48"),
   804 => (x"cc",x"7b",x"c0",x"87"),
   805 => (x"48",x"6e",x"49",x"a3"),
   806 => (x"66",x"c8",x"78",x"69"),
   807 => (x"cc",x"88",x"6b",x"48"),
   808 => (x"f0",x"c2",x"58",x"a6"),
   809 => (x"c8",x"48",x"bf",x"f0"),
   810 => (x"58",x"a6",x"c4",x"90"),
   811 => (x"6e",x"48",x"66",x"c8"),
   812 => (x"87",x"c9",x"01",x"a8"),
   813 => (x"6e",x"48",x"66",x"c8"),
   814 => (x"fd",x"c0",x"03",x"a8"),
   815 => (x"a3",x"c4",x"c1",x"87"),
   816 => (x"49",x"bf",x"6e",x"7e"),
   817 => (x"a1",x"75",x"91",x"c8"),
   818 => (x"79",x"66",x"cc",x"49"),
   819 => (x"c8",x"49",x"bf",x"6e"),
   820 => (x"49",x"a1",x"75",x"91"),
   821 => (x"79",x"66",x"81",x"c4"),
   822 => (x"6e",x"48",x"a6",x"d0"),
   823 => (x"66",x"d0",x"78",x"bf"),
   824 => (x"05",x"a8",x"c5",x"48"),
   825 => (x"a6",x"c4",x"87",x"c7"),
   826 => (x"c8",x"78",x"c0",x"48"),
   827 => (x"48",x"66",x"d0",x"87"),
   828 => (x"a6",x"c8",x"80",x"c1"),
   829 => (x"c4",x"48",x"6e",x"58"),
   830 => (x"66",x"c8",x"78",x"66"),
   831 => (x"f8",x"49",x"73",x"1e"),
   832 => (x"86",x"c4",x"87",x"ef"),
   833 => (x"1e",x"f0",x"e8",x"c2"),
   834 => (x"f1",x"f9",x"49",x"73"),
   835 => (x"49",x"a3",x"d0",x"87"),
   836 => (x"79",x"66",x"f0",x"c0"),
   837 => (x"4d",x"26",x"8e",x"e0"),
   838 => (x"4b",x"26",x"4c",x"26"),
   839 => (x"5e",x"0e",x"4f",x"26"),
   840 => (x"71",x"0e",x"5c",x"5b"),
   841 => (x"72",x"4b",x"c0",x"4a"),
   842 => (x"e0",x"c0",x"02",x"9a"),
   843 => (x"49",x"a2",x"da",x"87"),
   844 => (x"c2",x"4b",x"69",x"9f"),
   845 => (x"02",x"bf",x"f8",x"f0"),
   846 => (x"a2",x"d4",x"87",x"cf"),
   847 => (x"49",x"69",x"9f",x"49"),
   848 => (x"ff",x"ff",x"c0",x"4c"),
   849 => (x"c2",x"34",x"d0",x"9c"),
   850 => (x"74",x"4c",x"c0",x"87"),
   851 => (x"02",x"9b",x"73",x"b3"),
   852 => (x"c2",x"4a",x"87",x"df"),
   853 => (x"f0",x"f0",x"c2",x"8a"),
   854 => (x"c2",x"92",x"49",x"bf"),
   855 => (x"48",x"bf",x"d4",x"f5"),
   856 => (x"f5",x"c2",x"80",x"72"),
   857 => (x"48",x"71",x"58",x"f4"),
   858 => (x"f1",x"c2",x"30",x"c4"),
   859 => (x"e9",x"c0",x"58",x"c0"),
   860 => (x"d8",x"f5",x"c2",x"87"),
   861 => (x"f5",x"c2",x"4b",x"bf"),
   862 => (x"f5",x"c2",x"48",x"f0"),
   863 => (x"c2",x"78",x"bf",x"dc"),
   864 => (x"02",x"bf",x"f8",x"f0"),
   865 => (x"f0",x"c2",x"87",x"c9"),
   866 => (x"c4",x"49",x"bf",x"f0"),
   867 => (x"c2",x"87",x"c7",x"31"),
   868 => (x"49",x"bf",x"e0",x"f5"),
   869 => (x"f1",x"c2",x"31",x"c4"),
   870 => (x"f5",x"c2",x"59",x"c0"),
   871 => (x"4c",x"26",x"5b",x"f0"),
   872 => (x"4f",x"26",x"4b",x"26"),
   873 => (x"5c",x"5b",x"5e",x"0e"),
   874 => (x"86",x"f0",x"0e",x"5d"),
   875 => (x"cf",x"59",x"a6",x"c8"),
   876 => (x"f8",x"ff",x"ff",x"ff"),
   877 => (x"c4",x"7e",x"c0",x"4c"),
   878 => (x"87",x"d8",x"02",x"66"),
   879 => (x"48",x"ec",x"e8",x"c2"),
   880 => (x"e8",x"c2",x"78",x"c0"),
   881 => (x"f5",x"c2",x"48",x"e4"),
   882 => (x"c2",x"78",x"bf",x"f0"),
   883 => (x"c2",x"48",x"e8",x"e8"),
   884 => (x"78",x"bf",x"ec",x"f5"),
   885 => (x"48",x"cd",x"f1",x"c2"),
   886 => (x"f0",x"c2",x"50",x"c0"),
   887 => (x"c2",x"49",x"bf",x"fc"),
   888 => (x"4a",x"bf",x"ec",x"e8"),
   889 => (x"c4",x"03",x"aa",x"71"),
   890 => (x"49",x"72",x"87",x"cc"),
   891 => (x"c0",x"05",x"99",x"cf"),
   892 => (x"fe",x"c0",x"87",x"ea"),
   893 => (x"e8",x"c2",x"48",x"dc"),
   894 => (x"c2",x"78",x"bf",x"e4"),
   895 => (x"c2",x"1e",x"f0",x"e8"),
   896 => (x"49",x"bf",x"e4",x"e8"),
   897 => (x"48",x"e4",x"e8",x"c2"),
   898 => (x"71",x"78",x"a1",x"c1"),
   899 => (x"87",x"f2",x"df",x"ff"),
   900 => (x"fe",x"c0",x"86",x"c4"),
   901 => (x"e8",x"c2",x"48",x"d8"),
   902 => (x"87",x"cc",x"78",x"f0"),
   903 => (x"bf",x"d8",x"fe",x"c0"),
   904 => (x"80",x"e0",x"c0",x"48"),
   905 => (x"58",x"dc",x"fe",x"c0"),
   906 => (x"bf",x"ec",x"e8",x"c2"),
   907 => (x"c2",x"80",x"c1",x"48"),
   908 => (x"27",x"58",x"f0",x"e8"),
   909 => (x"00",x"00",x"0f",x"98"),
   910 => (x"4d",x"bf",x"97",x"bf"),
   911 => (x"e5",x"c2",x"02",x"9d"),
   912 => (x"ad",x"e5",x"c3",x"87"),
   913 => (x"87",x"de",x"c2",x"02"),
   914 => (x"bf",x"d8",x"fe",x"c0"),
   915 => (x"49",x"a3",x"cb",x"4b"),
   916 => (x"ac",x"cf",x"4c",x"11"),
   917 => (x"87",x"d2",x"c1",x"05"),
   918 => (x"99",x"df",x"49",x"75"),
   919 => (x"91",x"cd",x"89",x"c1"),
   920 => (x"81",x"c0",x"f1",x"c2"),
   921 => (x"12",x"4a",x"a3",x"c1"),
   922 => (x"4a",x"a3",x"c3",x"51"),
   923 => (x"a3",x"c5",x"51",x"12"),
   924 => (x"c7",x"51",x"12",x"4a"),
   925 => (x"51",x"12",x"4a",x"a3"),
   926 => (x"12",x"4a",x"a3",x"c9"),
   927 => (x"4a",x"a3",x"ce",x"51"),
   928 => (x"a3",x"d0",x"51",x"12"),
   929 => (x"d2",x"51",x"12",x"4a"),
   930 => (x"51",x"12",x"4a",x"a3"),
   931 => (x"12",x"4a",x"a3",x"d4"),
   932 => (x"4a",x"a3",x"d6",x"51"),
   933 => (x"a3",x"d8",x"51",x"12"),
   934 => (x"dc",x"51",x"12",x"4a"),
   935 => (x"51",x"12",x"4a",x"a3"),
   936 => (x"12",x"4a",x"a3",x"de"),
   937 => (x"c0",x"7e",x"c1",x"51"),
   938 => (x"49",x"74",x"87",x"fc"),
   939 => (x"c0",x"05",x"99",x"c8"),
   940 => (x"49",x"74",x"87",x"ed"),
   941 => (x"d3",x"05",x"99",x"d0"),
   942 => (x"66",x"e0",x"c0",x"87"),
   943 => (x"87",x"cc",x"c0",x"02"),
   944 => (x"e0",x"c0",x"49",x"73"),
   945 => (x"98",x"70",x"0f",x"66"),
   946 => (x"87",x"d3",x"c0",x"02"),
   947 => (x"c6",x"c0",x"05",x"6e"),
   948 => (x"c0",x"f1",x"c2",x"87"),
   949 => (x"c0",x"50",x"c0",x"48"),
   950 => (x"48",x"bf",x"d8",x"fe"),
   951 => (x"c2",x"87",x"e9",x"c2"),
   952 => (x"c0",x"48",x"cd",x"f1"),
   953 => (x"f0",x"c2",x"7e",x"50"),
   954 => (x"c2",x"49",x"bf",x"fc"),
   955 => (x"4a",x"bf",x"ec",x"e8"),
   956 => (x"fb",x"04",x"aa",x"71"),
   957 => (x"ff",x"cf",x"87",x"f4"),
   958 => (x"4c",x"f8",x"ff",x"ff"),
   959 => (x"bf",x"f0",x"f5",x"c2"),
   960 => (x"87",x"c8",x"c0",x"05"),
   961 => (x"bf",x"f8",x"f0",x"c2"),
   962 => (x"87",x"fa",x"c1",x"02"),
   963 => (x"bf",x"e8",x"e8",x"c2"),
   964 => (x"87",x"fd",x"ea",x"49"),
   965 => (x"58",x"ec",x"e8",x"c2"),
   966 => (x"c2",x"48",x"a6",x"c4"),
   967 => (x"78",x"bf",x"e8",x"e8"),
   968 => (x"bf",x"f8",x"f0",x"c2"),
   969 => (x"87",x"db",x"c0",x"02"),
   970 => (x"74",x"49",x"66",x"c4"),
   971 => (x"02",x"a9",x"74",x"99"),
   972 => (x"c8",x"87",x"c8",x"c0"),
   973 => (x"78",x"c0",x"48",x"a6"),
   974 => (x"c8",x"87",x"e7",x"c0"),
   975 => (x"78",x"c1",x"48",x"a6"),
   976 => (x"c4",x"87",x"df",x"c0"),
   977 => (x"ff",x"cf",x"49",x"66"),
   978 => (x"02",x"a9",x"99",x"f8"),
   979 => (x"cc",x"87",x"c8",x"c0"),
   980 => (x"78",x"c0",x"48",x"a6"),
   981 => (x"cc",x"87",x"c5",x"c0"),
   982 => (x"78",x"c1",x"48",x"a6"),
   983 => (x"cc",x"48",x"a6",x"c8"),
   984 => (x"66",x"c8",x"78",x"66"),
   985 => (x"87",x"de",x"c0",x"05"),
   986 => (x"c2",x"49",x"66",x"c4"),
   987 => (x"f0",x"f0",x"c2",x"89"),
   988 => (x"f5",x"c2",x"91",x"bf"),
   989 => (x"71",x"48",x"bf",x"d4"),
   990 => (x"e8",x"e8",x"c2",x"80"),
   991 => (x"ec",x"e8",x"c2",x"58"),
   992 => (x"f9",x"78",x"c0",x"48"),
   993 => (x"48",x"c0",x"87",x"d4"),
   994 => (x"ff",x"ff",x"ff",x"cf"),
   995 => (x"8e",x"f0",x"4c",x"f8"),
   996 => (x"4c",x"26",x"4d",x"26"),
   997 => (x"4f",x"26",x"4b",x"26"),
   998 => (x"00",x"00",x"00",x"00"),
   999 => (x"ff",x"ff",x"ff",x"ff"),
  1000 => (x"48",x"d4",x"ff",x"1e"),
  1001 => (x"68",x"78",x"ff",x"c3"),
  1002 => (x"1e",x"4f",x"26",x"48"),
  1003 => (x"c3",x"48",x"d4",x"ff"),
  1004 => (x"d0",x"ff",x"78",x"ff"),
  1005 => (x"78",x"e1",x"c0",x"48"),
  1006 => (x"d4",x"48",x"d4",x"ff"),
  1007 => (x"1e",x"4f",x"26",x"78"),
  1008 => (x"c0",x"48",x"d0",x"ff"),
  1009 => (x"4f",x"26",x"78",x"e0"),
  1010 => (x"87",x"d4",x"ff",x"1e"),
  1011 => (x"02",x"99",x"49",x"70"),
  1012 => (x"fb",x"c0",x"87",x"c6"),
  1013 => (x"87",x"f1",x"05",x"a9"),
  1014 => (x"4f",x"26",x"48",x"71"),
  1015 => (x"5c",x"5b",x"5e",x"0e"),
  1016 => (x"c0",x"4b",x"71",x"0e"),
  1017 => (x"87",x"f8",x"fe",x"4c"),
  1018 => (x"02",x"99",x"49",x"70"),
  1019 => (x"c0",x"87",x"f9",x"c0"),
  1020 => (x"c0",x"02",x"a9",x"ec"),
  1021 => (x"fb",x"c0",x"87",x"f2"),
  1022 => (x"eb",x"c0",x"02",x"a9"),
  1023 => (x"b7",x"66",x"cc",x"87"),
  1024 => (x"87",x"c7",x"03",x"ac"),
  1025 => (x"c2",x"02",x"66",x"d0"),
  1026 => (x"71",x"53",x"71",x"87"),
  1027 => (x"87",x"c2",x"02",x"99"),
  1028 => (x"cb",x"fe",x"84",x"c1"),
  1029 => (x"99",x"49",x"70",x"87"),
  1030 => (x"c0",x"87",x"cd",x"02"),
  1031 => (x"c7",x"02",x"a9",x"ec"),
  1032 => (x"a9",x"fb",x"c0",x"87"),
  1033 => (x"87",x"d5",x"ff",x"05"),
  1034 => (x"c3",x"02",x"66",x"d0"),
  1035 => (x"7b",x"97",x"c0",x"87"),
  1036 => (x"05",x"a9",x"fb",x"c0"),
  1037 => (x"4a",x"74",x"87",x"c7"),
  1038 => (x"c2",x"8a",x"0a",x"c0"),
  1039 => (x"72",x"4a",x"74",x"87"),
  1040 => (x"26",x"4c",x"26",x"48"),
  1041 => (x"1e",x"4f",x"26",x"4b"),
  1042 => (x"70",x"87",x"d5",x"fd"),
  1043 => (x"a9",x"f0",x"c0",x"49"),
  1044 => (x"c0",x"87",x"c9",x"04"),
  1045 => (x"c3",x"01",x"a9",x"f9"),
  1046 => (x"89",x"f0",x"c0",x"87"),
  1047 => (x"04",x"a9",x"c1",x"c1"),
  1048 => (x"da",x"c1",x"87",x"c9"),
  1049 => (x"87",x"c3",x"01",x"a9"),
  1050 => (x"71",x"89",x"f7",x"c0"),
  1051 => (x"0e",x"4f",x"26",x"48"),
  1052 => (x"5d",x"5c",x"5b",x"5e"),
  1053 => (x"71",x"86",x"f8",x"0e"),
  1054 => (x"fc",x"7e",x"c0",x"4c"),
  1055 => (x"4b",x"c0",x"87",x"ed"),
  1056 => (x"97",x"d0",x"c4",x"c1"),
  1057 => (x"a9",x"c0",x"49",x"bf"),
  1058 => (x"fc",x"87",x"cf",x"04"),
  1059 => (x"83",x"c1",x"87",x"fa"),
  1060 => (x"97",x"d0",x"c4",x"c1"),
  1061 => (x"06",x"ab",x"49",x"bf"),
  1062 => (x"c4",x"c1",x"87",x"f1"),
  1063 => (x"02",x"bf",x"97",x"d0"),
  1064 => (x"fb",x"fb",x"87",x"cf"),
  1065 => (x"99",x"49",x"70",x"87"),
  1066 => (x"c0",x"87",x"c6",x"02"),
  1067 => (x"f1",x"05",x"a9",x"ec"),
  1068 => (x"fb",x"4b",x"c0",x"87"),
  1069 => (x"4d",x"70",x"87",x"ea"),
  1070 => (x"c8",x"87",x"e5",x"fb"),
  1071 => (x"df",x"fb",x"58",x"a6"),
  1072 => (x"c1",x"4a",x"70",x"87"),
  1073 => (x"49",x"a4",x"c8",x"83"),
  1074 => (x"ad",x"49",x"69",x"97"),
  1075 => (x"c9",x"87",x"da",x"05"),
  1076 => (x"69",x"97",x"49",x"a4"),
  1077 => (x"a9",x"66",x"c4",x"49"),
  1078 => (x"ca",x"87",x"ce",x"05"),
  1079 => (x"69",x"97",x"49",x"a4"),
  1080 => (x"c4",x"05",x"aa",x"49"),
  1081 => (x"d0",x"7e",x"c1",x"87"),
  1082 => (x"ad",x"ec",x"c0",x"87"),
  1083 => (x"c0",x"87",x"c6",x"02"),
  1084 => (x"c4",x"05",x"ad",x"fb"),
  1085 => (x"c1",x"4b",x"c0",x"87"),
  1086 => (x"fe",x"02",x"6e",x"7e"),
  1087 => (x"fe",x"fa",x"87",x"f5"),
  1088 => (x"f8",x"48",x"73",x"87"),
  1089 => (x"26",x"4d",x"26",x"8e"),
  1090 => (x"26",x"4b",x"26",x"4c"),
  1091 => (x"00",x"00",x"00",x"4f"),
  1092 => (x"1e",x"73",x"1e",x"00"),
  1093 => (x"c8",x"4b",x"d4",x"ff"),
  1094 => (x"d0",x"ff",x"4a",x"66"),
  1095 => (x"78",x"c5",x"c8",x"48"),
  1096 => (x"c1",x"48",x"d4",x"ff"),
  1097 => (x"7b",x"11",x"78",x"d4"),
  1098 => (x"f9",x"05",x"8a",x"c1"),
  1099 => (x"48",x"d0",x"ff",x"87"),
  1100 => (x"4b",x"26",x"78",x"c4"),
  1101 => (x"5e",x"0e",x"4f",x"26"),
  1102 => (x"0e",x"5d",x"5c",x"5b"),
  1103 => (x"a6",x"c4",x"86",x"f8"),
  1104 => (x"c2",x"1e",x"6e",x"59"),
  1105 => (x"e3",x"49",x"c4",x"f6"),
  1106 => (x"86",x"c4",x"87",x"fe"),
  1107 => (x"c4",x"02",x"98",x"70"),
  1108 => (x"f2",x"c1",x"87",x"ee"),
  1109 => (x"6e",x"4c",x"bf",x"c8"),
  1110 => (x"87",x"d3",x"fc",x"49"),
  1111 => (x"c1",x"58",x"a6",x"c8"),
  1112 => (x"fe",x"1e",x"cc",x"ca"),
  1113 => (x"c4",x"87",x"e5",x"fc"),
  1114 => (x"c5",x"05",x"66",x"86"),
  1115 => (x"48",x"a6",x"c4",x"87"),
  1116 => (x"d0",x"ff",x"78",x"c1"),
  1117 => (x"ff",x"78",x"c5",x"48"),
  1118 => (x"d5",x"c1",x"48",x"d4"),
  1119 => (x"49",x"66",x"c4",x"78"),
  1120 => (x"31",x"c6",x"89",x"c1"),
  1121 => (x"97",x"c0",x"f2",x"c1"),
  1122 => (x"71",x"48",x"4a",x"bf"),
  1123 => (x"08",x"d4",x"ff",x"b0"),
  1124 => (x"48",x"d0",x"ff",x"78"),
  1125 => (x"f6",x"c2",x"78",x"c4"),
  1126 => (x"49",x"bf",x"97",x"c0"),
  1127 => (x"dd",x"02",x"99",x"d0"),
  1128 => (x"ff",x"78",x"c5",x"87"),
  1129 => (x"d6",x"c1",x"48",x"d4"),
  1130 => (x"ff",x"4a",x"c0",x"78"),
  1131 => (x"ff",x"c3",x"48",x"d4"),
  1132 => (x"c0",x"82",x"c1",x"78"),
  1133 => (x"f2",x"04",x"aa",x"e0"),
  1134 => (x"48",x"d0",x"ff",x"87"),
  1135 => (x"d4",x"ff",x"78",x"c4"),
  1136 => (x"78",x"ff",x"c3",x"48"),
  1137 => (x"c5",x"48",x"d0",x"ff"),
  1138 => (x"48",x"d4",x"ff",x"78"),
  1139 => (x"c1",x"78",x"d3",x"c1"),
  1140 => (x"48",x"d0",x"ff",x"78"),
  1141 => (x"b7",x"c0",x"78",x"c4"),
  1142 => (x"cc",x"c2",x"06",x"ac"),
  1143 => (x"cc",x"f6",x"c2",x"87"),
  1144 => (x"c4",x"8c",x"4b",x"bf"),
  1145 => (x"9b",x"73",x"5c",x"a6"),
  1146 => (x"87",x"dd",x"c1",x"02"),
  1147 => (x"8b",x"4d",x"c0",x"c8"),
  1148 => (x"03",x"ab",x"b7",x"c0"),
  1149 => (x"c0",x"c8",x"87",x"c6"),
  1150 => (x"4b",x"c0",x"4d",x"a3"),
  1151 => (x"97",x"c0",x"f6",x"c2"),
  1152 => (x"99",x"d0",x"49",x"bf"),
  1153 => (x"c0",x"87",x"cf",x"02"),
  1154 => (x"c4",x"f6",x"c2",x"1e"),
  1155 => (x"87",x"ee",x"e5",x"49"),
  1156 => (x"4c",x"70",x"86",x"c4"),
  1157 => (x"e8",x"c2",x"87",x"d8"),
  1158 => (x"f6",x"c2",x"1e",x"f0"),
  1159 => (x"dd",x"e5",x"49",x"c4"),
  1160 => (x"75",x"4c",x"70",x"87"),
  1161 => (x"f0",x"e8",x"c2",x"1e"),
  1162 => (x"87",x"e5",x"fb",x"49"),
  1163 => (x"9c",x"74",x"86",x"c8"),
  1164 => (x"c0",x"87",x"c5",x"05"),
  1165 => (x"87",x"ca",x"c1",x"48"),
  1166 => (x"f6",x"c2",x"1e",x"c1"),
  1167 => (x"f0",x"e3",x"49",x"c4"),
  1168 => (x"73",x"86",x"c4",x"87"),
  1169 => (x"e3",x"fe",x"05",x"9b"),
  1170 => (x"c0",x"4c",x"6e",x"87"),
  1171 => (x"d1",x"06",x"ac",x"b7"),
  1172 => (x"c4",x"f6",x"c2",x"87"),
  1173 => (x"d0",x"78",x"c0",x"48"),
  1174 => (x"f4",x"78",x"c0",x"80"),
  1175 => (x"d0",x"f6",x"c2",x"80"),
  1176 => (x"b7",x"c0",x"78",x"bf"),
  1177 => (x"f4",x"fd",x"01",x"ac"),
  1178 => (x"48",x"d0",x"ff",x"87"),
  1179 => (x"d4",x"ff",x"78",x"c5"),
  1180 => (x"78",x"d3",x"c1",x"48"),
  1181 => (x"d0",x"ff",x"78",x"c0"),
  1182 => (x"c1",x"78",x"c4",x"48"),
  1183 => (x"87",x"c2",x"c0",x"48"),
  1184 => (x"8e",x"f8",x"48",x"c0"),
  1185 => (x"4c",x"26",x"4d",x"26"),
  1186 => (x"4f",x"26",x"4b",x"26"),
  1187 => (x"20",x"74",x"6f",x"47"),
  1188 => (x"69",x"74",x"78",x"65"),
  1189 => (x"00",x"00",x"64",x"6e"),
  1190 => (x"64",x"61",x"6f",x"4c"),
  1191 => (x"2e",x"67",x"6e",x"69"),
  1192 => (x"00",x"00",x"2e",x"2e"),
  1193 => (x"61",x"42",x"20",x"80"),
  1194 => (x"00",x"00",x"6b",x"63"),
  1195 => (x"64",x"61",x"6f",x"4c"),
  1196 => (x"20",x"2e",x"2a",x"20"),
  1197 => (x"00",x"00",x"00",x"00"),
  1198 => (x"00",x"00",x"20",x"3a"),
  1199 => (x"61",x"42",x"20",x"80"),
  1200 => (x"00",x"00",x"6b",x"63"),
  1201 => (x"78",x"45",x"20",x"80"),
  1202 => (x"00",x"00",x"74",x"69"),
  1203 => (x"49",x"20",x"44",x"53"),
  1204 => (x"2e",x"74",x"69",x"6e"),
  1205 => (x"00",x"00",x"00",x"2e"),
  1206 => (x"00",x"00",x"4b",x"4f"),
  1207 => (x"54",x"4f",x"4f",x"42"),
  1208 => (x"20",x"20",x"20",x"20"),
  1209 => (x"00",x"4d",x"4f",x"52"),
  1210 => (x"5c",x"5b",x"5e",x"0e"),
  1211 => (x"86",x"fc",x"0e",x"5d"),
  1212 => (x"4b",x"c0",x"4d",x"71"),
  1213 => (x"c0",x"04",x"ad",x"4c"),
  1214 => (x"c1",x"c1",x"87",x"e8"),
  1215 => (x"9c",x"74",x"1e",x"ef"),
  1216 => (x"c0",x"87",x"c4",x"02"),
  1217 => (x"c1",x"87",x"c2",x"4a"),
  1218 => (x"ea",x"49",x"72",x"4a"),
  1219 => (x"86",x"c4",x"87",x"d6"),
  1220 => (x"83",x"c1",x"58",x"a6"),
  1221 => (x"87",x"c2",x"05",x"6e"),
  1222 => (x"84",x"c1",x"4b",x"75"),
  1223 => (x"ff",x"06",x"ab",x"75"),
  1224 => (x"48",x"6e",x"87",x"d8"),
  1225 => (x"4d",x"26",x"8e",x"fc"),
  1226 => (x"4b",x"26",x"4c",x"26"),
  1227 => (x"5e",x"0e",x"4f",x"26"),
  1228 => (x"71",x"0e",x"5c",x"5b"),
  1229 => (x"02",x"66",x"cc",x"4b"),
  1230 => (x"c0",x"4c",x"87",x"d8"),
  1231 => (x"d8",x"02",x"8c",x"f0"),
  1232 => (x"c1",x"4a",x"74",x"87"),
  1233 => (x"87",x"d1",x"02",x"8a"),
  1234 => (x"87",x"cd",x"02",x"8a"),
  1235 => (x"87",x"c9",x"02",x"8a"),
  1236 => (x"49",x"73",x"87",x"d9"),
  1237 => (x"d2",x"87",x"df",x"f7"),
  1238 => (x"c0",x"1e",x"74",x"87"),
  1239 => (x"f5",x"d7",x"c1",x"49"),
  1240 => (x"73",x"1e",x"74",x"87"),
  1241 => (x"ed",x"d7",x"c1",x"49"),
  1242 => (x"26",x"86",x"c8",x"87"),
  1243 => (x"26",x"4b",x"26",x"4c"),
  1244 => (x"5b",x"5e",x"0e",x"4f"),
  1245 => (x"fc",x"0e",x"5d",x"5c"),
  1246 => (x"49",x"4c",x"71",x"86"),
  1247 => (x"f7",x"c2",x"91",x"de"),
  1248 => (x"85",x"71",x"4d",x"e4"),
  1249 => (x"c1",x"02",x"6d",x"97"),
  1250 => (x"f7",x"c2",x"87",x"db"),
  1251 => (x"74",x"49",x"bf",x"d4"),
  1252 => (x"d3",x"fd",x"71",x"81"),
  1253 => (x"58",x"a6",x"c4",x"87"),
  1254 => (x"f2",x"c0",x"02",x"6e"),
  1255 => (x"d8",x"f7",x"c2",x"87"),
  1256 => (x"cb",x"4a",x"6e",x"4b"),
  1257 => (x"c3",x"fa",x"fe",x"49"),
  1258 => (x"cc",x"4b",x"74",x"87"),
  1259 => (x"cc",x"f2",x"c1",x"93"),
  1260 => (x"c1",x"83",x"c4",x"83"),
  1261 => (x"74",x"7b",x"d8",x"ca"),
  1262 => (x"db",x"c1",x"c1",x"49"),
  1263 => (x"c1",x"7b",x"75",x"87"),
  1264 => (x"bf",x"97",x"c4",x"f2"),
  1265 => (x"f7",x"c2",x"1e",x"49"),
  1266 => (x"e1",x"fd",x"49",x"d8"),
  1267 => (x"74",x"86",x"c4",x"87"),
  1268 => (x"c3",x"c1",x"c1",x"49"),
  1269 => (x"c1",x"49",x"c0",x"87"),
  1270 => (x"c2",x"87",x"df",x"c2"),
  1271 => (x"c0",x"48",x"fc",x"f5"),
  1272 => (x"ed",x"df",x"49",x"50"),
  1273 => (x"26",x"8e",x"fc",x"87"),
  1274 => (x"26",x"4c",x"26",x"4d"),
  1275 => (x"1e",x"4f",x"26",x"4b"),
  1276 => (x"4b",x"71",x"1e",x"73"),
  1277 => (x"d4",x"f7",x"c2",x"49"),
  1278 => (x"fb",x"71",x"81",x"bf"),
  1279 => (x"4a",x"70",x"87",x"ea"),
  1280 => (x"87",x"c4",x"02",x"9a"),
  1281 => (x"87",x"d6",x"e4",x"49"),
  1282 => (x"48",x"d4",x"f7",x"c2"),
  1283 => (x"49",x"73",x"78",x"c0"),
  1284 => (x"26",x"87",x"fa",x"c1"),
  1285 => (x"1e",x"4f",x"26",x"4b"),
  1286 => (x"4b",x"71",x"1e",x"73"),
  1287 => (x"02",x"4a",x"a3",x"c4"),
  1288 => (x"c1",x"87",x"d0",x"c1"),
  1289 => (x"87",x"dc",x"02",x"8a"),
  1290 => (x"f2",x"c0",x"02",x"8a"),
  1291 => (x"c1",x"05",x"8a",x"87"),
  1292 => (x"f7",x"c2",x"87",x"d3"),
  1293 => (x"c1",x"02",x"bf",x"d4"),
  1294 => (x"c1",x"48",x"87",x"cb"),
  1295 => (x"d8",x"f7",x"c2",x"88"),
  1296 => (x"87",x"c1",x"c1",x"58"),
  1297 => (x"bf",x"d4",x"f7",x"c2"),
  1298 => (x"c2",x"89",x"c6",x"49"),
  1299 => (x"c0",x"59",x"d8",x"f7"),
  1300 => (x"c0",x"03",x"a9",x"b7"),
  1301 => (x"f7",x"c2",x"87",x"ef"),
  1302 => (x"78",x"c0",x"48",x"d4"),
  1303 => (x"c2",x"87",x"e6",x"c0"),
  1304 => (x"02",x"bf",x"d0",x"f7"),
  1305 => (x"f7",x"c2",x"87",x"df"),
  1306 => (x"c1",x"48",x"bf",x"d4"),
  1307 => (x"d8",x"f7",x"c2",x"80"),
  1308 => (x"c2",x"87",x"d2",x"58"),
  1309 => (x"02",x"bf",x"d0",x"f7"),
  1310 => (x"f7",x"c2",x"87",x"cb"),
  1311 => (x"c6",x"48",x"bf",x"d4"),
  1312 => (x"d8",x"f7",x"c2",x"80"),
  1313 => (x"c4",x"49",x"73",x"58"),
  1314 => (x"26",x"4b",x"26",x"87"),
  1315 => (x"5b",x"5e",x"0e",x"4f"),
  1316 => (x"f0",x"0e",x"5d",x"5c"),
  1317 => (x"59",x"a6",x"d0",x"86"),
  1318 => (x"4d",x"f0",x"e8",x"c2"),
  1319 => (x"f7",x"c2",x"4c",x"c0"),
  1320 => (x"78",x"c1",x"48",x"d0"),
  1321 => (x"c0",x"48",x"a6",x"c8"),
  1322 => (x"5d",x"a6",x"c4",x"78"),
  1323 => (x"bf",x"d4",x"f7",x"c2"),
  1324 => (x"06",x"a8",x"c0",x"48"),
  1325 => (x"c8",x"87",x"c1",x"c1"),
  1326 => (x"a6",x"c4",x"5c",x"a6"),
  1327 => (x"f0",x"e8",x"c2",x"5d"),
  1328 => (x"c0",x"02",x"98",x"48"),
  1329 => (x"66",x"c4",x"87",x"f2"),
  1330 => (x"ef",x"c1",x"c1",x"4d"),
  1331 => (x"02",x"66",x"cc",x"1e"),
  1332 => (x"4c",x"c0",x"87",x"c4"),
  1333 => (x"4c",x"c1",x"87",x"c2"),
  1334 => (x"c7",x"e3",x"49",x"74"),
  1335 => (x"a6",x"86",x"c4",x"87"),
  1336 => (x"c8",x"85",x"c1",x"58"),
  1337 => (x"80",x"c1",x"48",x"66"),
  1338 => (x"c2",x"58",x"a6",x"cc"),
  1339 => (x"ad",x"bf",x"d4",x"f7"),
  1340 => (x"6e",x"87",x"c5",x"03"),
  1341 => (x"87",x"d1",x"ff",x"05"),
  1342 => (x"4c",x"c0",x"4d",x"6e"),
  1343 => (x"c3",x"02",x"9d",x"75"),
  1344 => (x"c1",x"c1",x"87",x"db"),
  1345 => (x"66",x"cc",x"1e",x"ef"),
  1346 => (x"c8",x"87",x"c7",x"02"),
  1347 => (x"78",x"c0",x"48",x"a6"),
  1348 => (x"a6",x"c8",x"87",x"c5"),
  1349 => (x"c8",x"78",x"c1",x"48"),
  1350 => (x"c7",x"e2",x"49",x"66"),
  1351 => (x"a6",x"86",x"c4",x"87"),
  1352 => (x"c2",x"02",x"6e",x"58"),
  1353 => (x"cb",x"49",x"87",x"e4"),
  1354 => (x"49",x"69",x"97",x"81"),
  1355 => (x"c1",x"02",x"99",x"d0"),
  1356 => (x"49",x"74",x"87",x"d4"),
  1357 => (x"f2",x"c1",x"91",x"cc"),
  1358 => (x"cf",x"c1",x"81",x"cc"),
  1359 => (x"81",x"c8",x"79",x"ef"),
  1360 => (x"74",x"51",x"ff",x"c3"),
  1361 => (x"c2",x"91",x"de",x"49"),
  1362 => (x"71",x"4d",x"e4",x"f7"),
  1363 => (x"97",x"c1",x"c2",x"85"),
  1364 => (x"49",x"a5",x"c1",x"7d"),
  1365 => (x"c2",x"51",x"e0",x"c0"),
  1366 => (x"bf",x"97",x"c0",x"f1"),
  1367 => (x"c1",x"87",x"d2",x"02"),
  1368 => (x"4b",x"a5",x"c2",x"84"),
  1369 => (x"4a",x"c0",x"f1",x"c2"),
  1370 => (x"f2",x"fe",x"49",x"db"),
  1371 => (x"d9",x"c1",x"87",x"fe"),
  1372 => (x"49",x"a5",x"cd",x"87"),
  1373 => (x"84",x"c1",x"51",x"c0"),
  1374 => (x"6e",x"4b",x"a5",x"c2"),
  1375 => (x"fe",x"49",x"cb",x"4a"),
  1376 => (x"c1",x"87",x"e9",x"f2"),
  1377 => (x"49",x"74",x"87",x"c4"),
  1378 => (x"f2",x"c1",x"91",x"cc"),
  1379 => (x"cd",x"c1",x"81",x"cc"),
  1380 => (x"f1",x"c2",x"79",x"f1"),
  1381 => (x"02",x"bf",x"97",x"c0"),
  1382 => (x"49",x"74",x"87",x"d8"),
  1383 => (x"84",x"c1",x"91",x"de"),
  1384 => (x"4b",x"e4",x"f7",x"c2"),
  1385 => (x"f1",x"c2",x"83",x"71"),
  1386 => (x"49",x"dd",x"4a",x"c0"),
  1387 => (x"87",x"fc",x"f1",x"fe"),
  1388 => (x"4b",x"74",x"87",x"d8"),
  1389 => (x"f7",x"c2",x"93",x"de"),
  1390 => (x"a3",x"cb",x"83",x"e4"),
  1391 => (x"c1",x"51",x"c0",x"49"),
  1392 => (x"4a",x"6e",x"73",x"84"),
  1393 => (x"f1",x"fe",x"49",x"cb"),
  1394 => (x"66",x"c8",x"87",x"e2"),
  1395 => (x"cc",x"80",x"c1",x"48"),
  1396 => (x"ac",x"c7",x"58",x"a6"),
  1397 => (x"87",x"c5",x"c0",x"03"),
  1398 => (x"e5",x"fc",x"05",x"6e"),
  1399 => (x"03",x"ac",x"c7",x"87"),
  1400 => (x"c2",x"87",x"e4",x"c0"),
  1401 => (x"c0",x"48",x"d0",x"f7"),
  1402 => (x"cc",x"49",x"74",x"78"),
  1403 => (x"cc",x"f2",x"c1",x"91"),
  1404 => (x"f1",x"cd",x"c1",x"81"),
  1405 => (x"de",x"49",x"74",x"79"),
  1406 => (x"e4",x"f7",x"c2",x"91"),
  1407 => (x"c1",x"51",x"c0",x"81"),
  1408 => (x"04",x"ac",x"c7",x"84"),
  1409 => (x"c1",x"87",x"dc",x"ff"),
  1410 => (x"c0",x"48",x"e8",x"f3"),
  1411 => (x"e0",x"f3",x"c1",x"50"),
  1412 => (x"ea",x"d9",x"c1",x"48"),
  1413 => (x"c1",x"80",x"c4",x"78"),
  1414 => (x"c8",x"78",x"e4",x"ca"),
  1415 => (x"d7",x"d0",x"c1",x"80"),
  1416 => (x"49",x"66",x"cc",x"78"),
  1417 => (x"87",x"f0",x"f7",x"c0"),
  1418 => (x"4d",x"26",x"8e",x"f0"),
  1419 => (x"4b",x"26",x"4c",x"26"),
  1420 => (x"73",x"1e",x"4f",x"26"),
  1421 => (x"49",x"4b",x"71",x"1e"),
  1422 => (x"f2",x"c1",x"91",x"cc"),
  1423 => (x"a1",x"c8",x"81",x"cc"),
  1424 => (x"c0",x"f2",x"c1",x"4a"),
  1425 => (x"c9",x"50",x"12",x"48"),
  1426 => (x"c4",x"c1",x"4a",x"a1"),
  1427 => (x"50",x"12",x"48",x"d0"),
  1428 => (x"f2",x"c1",x"81",x"ca"),
  1429 => (x"50",x"11",x"48",x"c4"),
  1430 => (x"f0",x"f8",x"49",x"73"),
  1431 => (x"26",x"4b",x"26",x"87"),
  1432 => (x"49",x"c0",x"1e",x"4f"),
  1433 => (x"87",x"d2",x"f8",x"c0"),
  1434 => (x"71",x"1e",x"4f",x"26"),
  1435 => (x"91",x"cc",x"49",x"4a"),
  1436 => (x"81",x"cc",x"f2",x"c1"),
  1437 => (x"f5",x"c2",x"81",x"c8"),
  1438 => (x"50",x"11",x"48",x"fc"),
  1439 => (x"49",x"a2",x"f0",x"c0"),
  1440 => (x"87",x"f3",x"ec",x"fe"),
  1441 => (x"c9",x"d5",x"49",x"c0"),
  1442 => (x"1e",x"4f",x"26",x"87"),
  1443 => (x"c3",x"4a",x"d4",x"ff"),
  1444 => (x"d0",x"ff",x"7a",x"ff"),
  1445 => (x"78",x"e1",x"c0",x"48"),
  1446 => (x"7a",x"71",x"7a",x"de"),
  1447 => (x"28",x"b7",x"c8",x"48"),
  1448 => (x"48",x"71",x"7a",x"70"),
  1449 => (x"70",x"28",x"b7",x"d0"),
  1450 => (x"d8",x"48",x"71",x"7a"),
  1451 => (x"7a",x"70",x"28",x"b7"),
  1452 => (x"c0",x"48",x"d0",x"ff"),
  1453 => (x"4f",x"26",x"78",x"e0"),
  1454 => (x"5c",x"5b",x"5e",x"0e"),
  1455 => (x"86",x"f4",x"0e",x"5d"),
  1456 => (x"cc",x"49",x"4d",x"71"),
  1457 => (x"cc",x"f2",x"c1",x"91"),
  1458 => (x"4a",x"a1",x"c8",x"81"),
  1459 => (x"c4",x"7e",x"a1",x"ca"),
  1460 => (x"f5",x"c2",x"48",x"a6"),
  1461 => (x"6e",x"78",x"bf",x"f8"),
  1462 => (x"c4",x"4b",x"bf",x"97"),
  1463 => (x"2c",x"73",x"4c",x"66"),
  1464 => (x"a6",x"cc",x"48",x"12"),
  1465 => (x"c1",x"9c",x"70",x"58"),
  1466 => (x"97",x"81",x"c9",x"84"),
  1467 => (x"ac",x"b7",x"49",x"69"),
  1468 => (x"c0",x"87",x"c2",x"04"),
  1469 => (x"bf",x"97",x"6e",x"4c"),
  1470 => (x"49",x"66",x"c8",x"4a"),
  1471 => (x"b9",x"ff",x"31",x"72"),
  1472 => (x"74",x"99",x"66",x"c4"),
  1473 => (x"70",x"30",x"72",x"48"),
  1474 => (x"f5",x"c2",x"b1",x"4a"),
  1475 => (x"fd",x"71",x"59",x"fc"),
  1476 => (x"1e",x"c7",x"87",x"f9"),
  1477 => (x"bf",x"cc",x"f7",x"c2"),
  1478 => (x"cc",x"f2",x"c1",x"1e"),
  1479 => (x"fc",x"f5",x"c2",x"1e"),
  1480 => (x"c1",x"49",x"bf",x"97"),
  1481 => (x"49",x"75",x"87",x"f4"),
  1482 => (x"87",x"ec",x"f3",x"c0"),
  1483 => (x"4d",x"26",x"8e",x"e8"),
  1484 => (x"4b",x"26",x"4c",x"26"),
  1485 => (x"73",x"1e",x"4f",x"26"),
  1486 => (x"49",x"4b",x"71",x"1e"),
  1487 => (x"73",x"87",x"f9",x"fd"),
  1488 => (x"87",x"f4",x"fd",x"49"),
  1489 => (x"4f",x"26",x"4b",x"26"),
  1490 => (x"71",x"1e",x"73",x"1e"),
  1491 => (x"4a",x"a3",x"c2",x"4b"),
  1492 => (x"c1",x"87",x"d6",x"02"),
  1493 => (x"e2",x"c0",x"05",x"8a"),
  1494 => (x"cc",x"f7",x"c2",x"87"),
  1495 => (x"87",x"db",x"02",x"bf"),
  1496 => (x"c2",x"88",x"c1",x"48"),
  1497 => (x"d2",x"58",x"d0",x"f7"),
  1498 => (x"d0",x"f7",x"c2",x"87"),
  1499 => (x"87",x"cb",x"02",x"bf"),
  1500 => (x"bf",x"cc",x"f7",x"c2"),
  1501 => (x"c2",x"80",x"c1",x"48"),
  1502 => (x"c7",x"58",x"d0",x"f7"),
  1503 => (x"cc",x"f7",x"c2",x"1e"),
  1504 => (x"f2",x"c1",x"1e",x"bf"),
  1505 => (x"f5",x"c2",x"1e",x"cc"),
  1506 => (x"49",x"bf",x"97",x"fc"),
  1507 => (x"49",x"73",x"87",x"cc"),
  1508 => (x"87",x"c4",x"f2",x"c0"),
  1509 => (x"4b",x"26",x"8e",x"f4"),
  1510 => (x"5e",x"0e",x"4f",x"26"),
  1511 => (x"0e",x"5d",x"5c",x"5b"),
  1512 => (x"c0",x"86",x"cc",x"ff"),
  1513 => (x"cc",x"59",x"a6",x"e8"),
  1514 => (x"78",x"c0",x"48",x"a6"),
  1515 => (x"78",x"c0",x"80",x"c4"),
  1516 => (x"78",x"c0",x"80",x"c4"),
  1517 => (x"c8",x"c1",x"80",x"c4"),
  1518 => (x"80",x"c4",x"78",x"66"),
  1519 => (x"80",x"c4",x"78",x"c1"),
  1520 => (x"f7",x"c2",x"78",x"c1"),
  1521 => (x"78",x"c1",x"48",x"d0"),
  1522 => (x"87",x"df",x"df",x"ff"),
  1523 => (x"87",x"f8",x"df",x"ff"),
  1524 => (x"87",x"cc",x"df",x"ff"),
  1525 => (x"fb",x"c0",x"4d",x"70"),
  1526 => (x"f3",x"c1",x"02",x"ad"),
  1527 => (x"66",x"e4",x"c0",x"87"),
  1528 => (x"87",x"e8",x"c1",x"05"),
  1529 => (x"4a",x"66",x"c4",x"c1"),
  1530 => (x"7e",x"6a",x"82",x"c4"),
  1531 => (x"48",x"ec",x"ca",x"c1"),
  1532 => (x"41",x"20",x"49",x"6e"),
  1533 => (x"51",x"10",x"41",x"20"),
  1534 => (x"48",x"66",x"c4",x"c1"),
  1535 => (x"78",x"f2",x"d8",x"c1"),
  1536 => (x"81",x"c7",x"49",x"6a"),
  1537 => (x"c4",x"c1",x"51",x"75"),
  1538 => (x"81",x"c8",x"49",x"66"),
  1539 => (x"a6",x"dc",x"51",x"c1"),
  1540 => (x"c1",x"78",x"c2",x"48"),
  1541 => (x"c9",x"49",x"66",x"c4"),
  1542 => (x"c1",x"51",x"c0",x"81"),
  1543 => (x"ca",x"49",x"66",x"c4"),
  1544 => (x"c1",x"51",x"c0",x"81"),
  1545 => (x"6a",x"1e",x"d8",x"1e"),
  1546 => (x"ff",x"81",x"c8",x"49"),
  1547 => (x"c8",x"87",x"ed",x"de"),
  1548 => (x"66",x"c8",x"c1",x"86"),
  1549 => (x"01",x"a8",x"c0",x"48"),
  1550 => (x"a6",x"d4",x"87",x"c7"),
  1551 => (x"cf",x"78",x"c1",x"48"),
  1552 => (x"66",x"c8",x"c1",x"87"),
  1553 => (x"dc",x"88",x"c1",x"48"),
  1554 => (x"87",x"c4",x"58",x"a6"),
  1555 => (x"87",x"f8",x"dd",x"ff"),
  1556 => (x"cb",x"02",x"9d",x"75"),
  1557 => (x"66",x"d4",x"87",x"f6"),
  1558 => (x"66",x"cc",x"c1",x"48"),
  1559 => (x"eb",x"cb",x"03",x"a8"),
  1560 => (x"ff",x"7e",x"c0",x"87"),
  1561 => (x"70",x"87",x"f9",x"dc"),
  1562 => (x"c6",x"c1",x"48",x"4d"),
  1563 => (x"58",x"a6",x"c8",x"88"),
  1564 => (x"c1",x"02",x"98",x"70"),
  1565 => (x"c9",x"48",x"87",x"d7"),
  1566 => (x"58",x"a6",x"c8",x"88"),
  1567 => (x"c5",x"02",x"98",x"70"),
  1568 => (x"c1",x"48",x"87",x"da"),
  1569 => (x"58",x"a6",x"c8",x"88"),
  1570 => (x"c2",x"02",x"98",x"70"),
  1571 => (x"c3",x"48",x"87",x"f9"),
  1572 => (x"58",x"a6",x"c8",x"88"),
  1573 => (x"cf",x"02",x"98",x"70"),
  1574 => (x"88",x"c1",x"48",x"87"),
  1575 => (x"70",x"58",x"a6",x"c8"),
  1576 => (x"f7",x"c4",x"02",x"98"),
  1577 => (x"87",x"c3",x"ca",x"87"),
  1578 => (x"ff",x"7e",x"f0",x"c0"),
  1579 => (x"70",x"87",x"f1",x"db"),
  1580 => (x"ad",x"ec",x"c0",x"4d"),
  1581 => (x"c4",x"87",x"c3",x"02"),
  1582 => (x"ec",x"c0",x"5d",x"a6"),
  1583 => (x"87",x"cd",x"02",x"ad"),
  1584 => (x"87",x"dc",x"db",x"ff"),
  1585 => (x"ec",x"c0",x"4d",x"70"),
  1586 => (x"f3",x"ff",x"05",x"ad"),
  1587 => (x"66",x"e4",x"c0",x"87"),
  1588 => (x"87",x"ea",x"c1",x"05"),
  1589 => (x"02",x"ad",x"ec",x"c0"),
  1590 => (x"db",x"ff",x"87",x"c4"),
  1591 => (x"1e",x"c0",x"87",x"c2"),
  1592 => (x"66",x"dc",x"1e",x"ca"),
  1593 => (x"c1",x"93",x"cc",x"4b"),
  1594 => (x"c4",x"83",x"66",x"cc"),
  1595 => (x"49",x"6c",x"4c",x"a3"),
  1596 => (x"87",x"e8",x"db",x"ff"),
  1597 => (x"1e",x"de",x"1e",x"c1"),
  1598 => (x"db",x"ff",x"49",x"6c"),
  1599 => (x"86",x"d0",x"87",x"de"),
  1600 => (x"7b",x"f2",x"d8",x"c1"),
  1601 => (x"dc",x"49",x"a3",x"c8"),
  1602 => (x"a3",x"c9",x"51",x"66"),
  1603 => (x"66",x"e0",x"c0",x"49"),
  1604 => (x"49",x"a3",x"ca",x"51"),
  1605 => (x"66",x"dc",x"51",x"6e"),
  1606 => (x"c0",x"80",x"c1",x"48"),
  1607 => (x"d4",x"58",x"a6",x"e0"),
  1608 => (x"66",x"d8",x"48",x"66"),
  1609 => (x"87",x"cb",x"04",x"a8"),
  1610 => (x"c1",x"48",x"66",x"d4"),
  1611 => (x"58",x"a6",x"d8",x"80"),
  1612 => (x"d8",x"87",x"fe",x"c7"),
  1613 => (x"88",x"c1",x"48",x"66"),
  1614 => (x"c7",x"58",x"a6",x"dc"),
  1615 => (x"da",x"ff",x"87",x"f3"),
  1616 => (x"4d",x"70",x"87",x"c6"),
  1617 => (x"ff",x"87",x"ea",x"c7"),
  1618 => (x"d0",x"87",x"fc",x"db"),
  1619 => (x"66",x"d0",x"58",x"a6"),
  1620 => (x"c6",x"c0",x"06",x"a8"),
  1621 => (x"48",x"a6",x"d0",x"87"),
  1622 => (x"ff",x"78",x"66",x"cc"),
  1623 => (x"c0",x"87",x"e8",x"db"),
  1624 => (x"c1",x"05",x"a8",x"ec"),
  1625 => (x"e4",x"c0",x"87",x"f6"),
  1626 => (x"e6",x"c1",x"05",x"66"),
  1627 => (x"49",x"66",x"d4",x"87"),
  1628 => (x"c4",x"c1",x"91",x"cc"),
  1629 => (x"a1",x"c4",x"81",x"66"),
  1630 => (x"c8",x"4c",x"6a",x"4a"),
  1631 => (x"66",x"cc",x"4a",x"a1"),
  1632 => (x"ea",x"d9",x"c1",x"52"),
  1633 => (x"d7",x"d8",x"ff",x"79"),
  1634 => (x"9d",x"4d",x"70",x"87"),
  1635 => (x"c0",x"87",x"db",x"02"),
  1636 => (x"c0",x"02",x"ad",x"fb"),
  1637 => (x"54",x"75",x"87",x"d4"),
  1638 => (x"87",x"c4",x"d8",x"ff"),
  1639 => (x"02",x"9d",x"4d",x"70"),
  1640 => (x"c0",x"87",x"c7",x"c0"),
  1641 => (x"ff",x"05",x"ad",x"fb"),
  1642 => (x"e0",x"c0",x"87",x"ec"),
  1643 => (x"54",x"c1",x"c2",x"54"),
  1644 => (x"d4",x"7c",x"97",x"c0"),
  1645 => (x"66",x"d8",x"48",x"66"),
  1646 => (x"cb",x"c0",x"04",x"a8"),
  1647 => (x"48",x"66",x"d4",x"87"),
  1648 => (x"a6",x"d8",x"80",x"c1"),
  1649 => (x"87",x"e9",x"c5",x"58"),
  1650 => (x"c1",x"48",x"66",x"d8"),
  1651 => (x"58",x"a6",x"dc",x"88"),
  1652 => (x"ff",x"87",x"de",x"c5"),
  1653 => (x"70",x"87",x"f1",x"d7"),
  1654 => (x"87",x"d5",x"c5",x"4d"),
  1655 => (x"c0",x"48",x"66",x"cc"),
  1656 => (x"05",x"a8",x"66",x"e4"),
  1657 => (x"c0",x"87",x"f6",x"c4"),
  1658 => (x"c0",x"48",x"a6",x"e8"),
  1659 => (x"d6",x"d9",x"ff",x"78"),
  1660 => (x"58",x"a6",x"c4",x"87"),
  1661 => (x"87",x"cf",x"d9",x"ff"),
  1662 => (x"58",x"a6",x"f0",x"c0"),
  1663 => (x"05",x"a8",x"ec",x"c0"),
  1664 => (x"a6",x"87",x"c7",x"c0"),
  1665 => (x"c0",x"78",x"6e",x"48"),
  1666 => (x"d6",x"ff",x"87",x"c4"),
  1667 => (x"66",x"d4",x"87",x"d2"),
  1668 => (x"c1",x"91",x"cc",x"49"),
  1669 => (x"71",x"48",x"66",x"c4"),
  1670 => (x"58",x"a6",x"c8",x"80"),
  1671 => (x"c8",x"4a",x"66",x"c4"),
  1672 => (x"49",x"66",x"c4",x"82"),
  1673 => (x"51",x"6e",x"81",x"ca"),
  1674 => (x"49",x"66",x"ec",x"c0"),
  1675 => (x"89",x"6e",x"81",x"c1"),
  1676 => (x"30",x"71",x"48",x"c1"),
  1677 => (x"89",x"c1",x"49",x"70"),
  1678 => (x"c2",x"7a",x"97",x"71"),
  1679 => (x"49",x"bf",x"f8",x"f5"),
  1680 => (x"6a",x"97",x"29",x"6e"),
  1681 => (x"98",x"71",x"48",x"4a"),
  1682 => (x"58",x"a6",x"f4",x"c0"),
  1683 => (x"c4",x"48",x"66",x"c4"),
  1684 => (x"58",x"a6",x"cc",x"80"),
  1685 => (x"4c",x"bf",x"66",x"c8"),
  1686 => (x"48",x"66",x"e4",x"c0"),
  1687 => (x"02",x"a8",x"66",x"cc"),
  1688 => (x"c0",x"87",x"c5",x"c0"),
  1689 => (x"87",x"c2",x"c0",x"7e"),
  1690 => (x"1e",x"6e",x"7e",x"c1"),
  1691 => (x"74",x"1e",x"e0",x"c0"),
  1692 => (x"e7",x"d5",x"ff",x"49"),
  1693 => (x"70",x"86",x"c8",x"87"),
  1694 => (x"ad",x"b7",x"c0",x"4d"),
  1695 => (x"87",x"d5",x"c1",x"06"),
  1696 => (x"66",x"c8",x"84",x"75"),
  1697 => (x"e0",x"c0",x"49",x"bf"),
  1698 => (x"4b",x"89",x"74",x"81"),
  1699 => (x"4a",x"f8",x"ca",x"c1"),
  1700 => (x"d7",x"de",x"fe",x"71"),
  1701 => (x"c4",x"84",x"c2",x"87"),
  1702 => (x"e8",x"c0",x"5c",x"a6"),
  1703 => (x"80",x"c1",x"48",x"66"),
  1704 => (x"58",x"a6",x"ec",x"c0"),
  1705 => (x"49",x"66",x"f0",x"c0"),
  1706 => (x"a9",x"70",x"81",x"c1"),
  1707 => (x"87",x"c5",x"c0",x"02"),
  1708 => (x"c2",x"c0",x"4c",x"c0"),
  1709 => (x"74",x"4c",x"c1",x"87"),
  1710 => (x"bf",x"66",x"cc",x"1e"),
  1711 => (x"81",x"e0",x"c0",x"49"),
  1712 => (x"71",x"89",x"66",x"c4"),
  1713 => (x"49",x"66",x"c8",x"1e"),
  1714 => (x"87",x"d0",x"d4",x"ff"),
  1715 => (x"b7",x"c0",x"86",x"c8"),
  1716 => (x"c5",x"ff",x"01",x"a8"),
  1717 => (x"66",x"e8",x"c0",x"87"),
  1718 => (x"87",x"d3",x"c0",x"02"),
  1719 => (x"c9",x"49",x"66",x"c4"),
  1720 => (x"66",x"e8",x"c0",x"81"),
  1721 => (x"48",x"66",x"c4",x"51"),
  1722 => (x"78",x"f8",x"da",x"c1"),
  1723 => (x"c4",x"87",x"ce",x"c0"),
  1724 => (x"81",x"c9",x"49",x"66"),
  1725 => (x"66",x"c4",x"51",x"c2"),
  1726 => (x"f6",x"dc",x"c1",x"48"),
  1727 => (x"48",x"66",x"d4",x"78"),
  1728 => (x"04",x"a8",x"66",x"d8"),
  1729 => (x"d4",x"87",x"cb",x"c0"),
  1730 => (x"80",x"c1",x"48",x"66"),
  1731 => (x"c0",x"58",x"a6",x"d8"),
  1732 => (x"66",x"d8",x"87",x"d1"),
  1733 => (x"dc",x"88",x"c1",x"48"),
  1734 => (x"c6",x"c0",x"58",x"a6"),
  1735 => (x"e7",x"d2",x"ff",x"87"),
  1736 => (x"cc",x"4d",x"70",x"87"),
  1737 => (x"78",x"c0",x"48",x"a6"),
  1738 => (x"ff",x"87",x"c6",x"c0"),
  1739 => (x"70",x"87",x"d9",x"d2"),
  1740 => (x"66",x"e0",x"c0",x"4d"),
  1741 => (x"c0",x"80",x"c1",x"48"),
  1742 => (x"75",x"58",x"a6",x"e4"),
  1743 => (x"cb",x"c0",x"02",x"9d"),
  1744 => (x"48",x"66",x"d4",x"87"),
  1745 => (x"a8",x"66",x"cc",x"c1"),
  1746 => (x"87",x"d5",x"f4",x"04"),
  1747 => (x"c7",x"48",x"66",x"d4"),
  1748 => (x"e1",x"c0",x"03",x"a8"),
  1749 => (x"4c",x"66",x"d4",x"87"),
  1750 => (x"48",x"d0",x"f7",x"c2"),
  1751 => (x"49",x"74",x"78",x"c0"),
  1752 => (x"c4",x"c1",x"91",x"cc"),
  1753 => (x"a1",x"c4",x"81",x"66"),
  1754 => (x"c0",x"4a",x"6a",x"4a"),
  1755 => (x"84",x"c1",x"79",x"52"),
  1756 => (x"ff",x"04",x"ac",x"c7"),
  1757 => (x"e4",x"c0",x"87",x"e2"),
  1758 => (x"e2",x"c0",x"02",x"66"),
  1759 => (x"66",x"c4",x"c1",x"87"),
  1760 => (x"81",x"d4",x"c1",x"49"),
  1761 => (x"4a",x"66",x"c4",x"c1"),
  1762 => (x"c0",x"82",x"dc",x"c1"),
  1763 => (x"ea",x"d9",x"c1",x"52"),
  1764 => (x"66",x"c4",x"c1",x"79"),
  1765 => (x"81",x"d8",x"c1",x"49"),
  1766 => (x"79",x"fc",x"ca",x"c1"),
  1767 => (x"c1",x"87",x"d6",x"c0"),
  1768 => (x"c1",x"49",x"66",x"c4"),
  1769 => (x"c4",x"c1",x"81",x"d4"),
  1770 => (x"d8",x"c1",x"4a",x"66"),
  1771 => (x"c4",x"cb",x"c1",x"82"),
  1772 => (x"e1",x"d9",x"c1",x"7a"),
  1773 => (x"66",x"c4",x"c1",x"79"),
  1774 => (x"81",x"e0",x"c1",x"49"),
  1775 => (x"79",x"c8",x"dd",x"c1"),
  1776 => (x"87",x"fb",x"cf",x"ff"),
  1777 => (x"ff",x"48",x"66",x"d0"),
  1778 => (x"4d",x"26",x"8e",x"cc"),
  1779 => (x"4b",x"26",x"4c",x"26"),
  1780 => (x"c7",x"1e",x"4f",x"26"),
  1781 => (x"cc",x"f7",x"c2",x"1e"),
  1782 => (x"f2",x"c1",x"1e",x"bf"),
  1783 => (x"f5",x"c2",x"1e",x"cc"),
  1784 => (x"49",x"bf",x"97",x"fc"),
  1785 => (x"c1",x"87",x"f3",x"ee"),
  1786 => (x"c0",x"49",x"cc",x"f2"),
  1787 => (x"f4",x"87",x"f8",x"e1"),
  1788 => (x"1e",x"4f",x"26",x"8e"),
  1789 => (x"48",x"c0",x"f2",x"c1"),
  1790 => (x"f3",x"c1",x"50",x"c0"),
  1791 => (x"ff",x"49",x"bf",x"f8"),
  1792 => (x"c0",x"87",x"f3",x"d4"),
  1793 => (x"1e",x"4f",x"26",x"48"),
  1794 => (x"d4",x"c7",x"1e",x"73"),
  1795 => (x"d8",x"f7",x"c2",x"87"),
  1796 => (x"ff",x"50",x"c0",x"48"),
  1797 => (x"ff",x"c3",x"48",x"d4"),
  1798 => (x"cc",x"cb",x"c1",x"78"),
  1799 => (x"f2",x"d6",x"fe",x"49"),
  1800 => (x"c7",x"e2",x"fe",x"87"),
  1801 => (x"02",x"98",x"70",x"87"),
  1802 => (x"eb",x"fe",x"87",x"cd"),
  1803 => (x"98",x"70",x"87",x"e5"),
  1804 => (x"c1",x"87",x"c4",x"02"),
  1805 => (x"c0",x"87",x"c2",x"4a"),
  1806 => (x"02",x"9a",x"72",x"4a"),
  1807 => (x"cb",x"c1",x"87",x"c8"),
  1808 => (x"d6",x"fe",x"49",x"d8"),
  1809 => (x"f7",x"c2",x"87",x"cd"),
  1810 => (x"78",x"c0",x"48",x"cc"),
  1811 => (x"48",x"fc",x"f5",x"c2"),
  1812 => (x"fd",x"49",x"50",x"c0"),
  1813 => (x"da",x"fe",x"87",x"fc"),
  1814 => (x"9b",x"4b",x"70",x"87"),
  1815 => (x"c1",x"87",x"cf",x"02"),
  1816 => (x"c7",x"5b",x"e8",x"f3"),
  1817 => (x"87",x"f0",x"de",x"49"),
  1818 => (x"e0",x"c0",x"49",x"c1"),
  1819 => (x"f3",x"c2",x"87",x"cc"),
  1820 => (x"d2",x"e1",x"c0",x"87"),
  1821 => (x"eb",x"ef",x"c0",x"87"),
  1822 => (x"87",x"f5",x"ff",x"87"),
  1823 => (x"4f",x"26",x"4b",x"26"),
  1824 => (x"00",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"00",x"00"),
  1826 => (x"00",x"00",x"00",x"01"),
  1827 => (x"00",x"00",x"13",x"71"),
  1828 => (x"00",x"00",x"2d",x"e4"),
  1829 => (x"d4",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"13",x"71"),
  1831 => (x"00",x"00",x"2e",x"02"),
  1832 => (x"d4",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"13",x"71"),
  1834 => (x"00",x"00",x"2e",x"20"),
  1835 => (x"d4",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"13",x"71"),
  1837 => (x"00",x"00",x"2e",x"3e"),
  1838 => (x"d4",x"00",x"00",x"00"),
  1839 => (x"00",x"00",x"13",x"71"),
  1840 => (x"00",x"00",x"2e",x"5c"),
  1841 => (x"d4",x"00",x"00",x"00"),
  1842 => (x"00",x"00",x"13",x"71"),
  1843 => (x"00",x"00",x"2e",x"7a"),
  1844 => (x"d4",x"00",x"00",x"00"),
  1845 => (x"00",x"00",x"13",x"71"),
  1846 => (x"00",x"00",x"2e",x"98"),
  1847 => (x"d4",x"00",x"00",x"00"),
  1848 => (x"00",x"00",x"16",x"6a"),
  1849 => (x"00",x"00",x"00",x"00"),
  1850 => (x"d4",x"00",x"00",x"00"),
  1851 => (x"00",x"00",x"14",x"17"),
  1852 => (x"00",x"00",x"00",x"00"),
  1853 => (x"d4",x"00",x"00",x"00"),
  1854 => (x"00",x"00",x"12",x"dc"),
  1855 => (x"dc",x"86",x"fc",x"1e"),
  1856 => (x"58",x"a6",x"c4",x"87"),
  1857 => (x"4f",x"26",x"8e",x"fc"),
  1858 => (x"48",x"f0",x"fe",x"1e"),
  1859 => (x"09",x"cd",x"78",x"c0"),
  1860 => (x"4f",x"26",x"09",x"79"),
  1861 => (x"fc",x"f3",x"c1",x"1e"),
  1862 => (x"26",x"87",x"ed",x"49"),
  1863 => (x"f0",x"fe",x"1e",x"4f"),
  1864 => (x"4f",x"26",x"48",x"bf"),
  1865 => (x"48",x"f0",x"fe",x"1e"),
  1866 => (x"4f",x"26",x"78",x"c1"),
  1867 => (x"48",x"f0",x"fe",x"1e"),
  1868 => (x"4f",x"26",x"78",x"c0"),
  1869 => (x"c0",x"4a",x"71",x"1e"),
  1870 => (x"4f",x"26",x"51",x"52"),
  1871 => (x"5c",x"5b",x"5e",x"0e"),
  1872 => (x"86",x"f4",x"0e",x"5d"),
  1873 => (x"6d",x"97",x"4d",x"71"),
  1874 => (x"58",x"a6",x"c4",x"48"),
  1875 => (x"97",x"4c",x"a5",x"c1"),
  1876 => (x"a6",x"c8",x"48",x"6c"),
  1877 => (x"c4",x"48",x"6e",x"58"),
  1878 => (x"c5",x"05",x"a8",x"66"),
  1879 => (x"c0",x"48",x"ff",x"87"),
  1880 => (x"c7",x"ff",x"87",x"e7"),
  1881 => (x"49",x"a5",x"c2",x"87"),
  1882 => (x"71",x"4b",x"6c",x"97"),
  1883 => (x"6b",x"97",x"4b",x"a3"),
  1884 => (x"48",x"6c",x"97",x"4b"),
  1885 => (x"c1",x"58",x"a6",x"c4"),
  1886 => (x"58",x"a6",x"c8",x"80"),
  1887 => (x"a6",x"cc",x"98",x"c7"),
  1888 => (x"7c",x"97",x"70",x"58"),
  1889 => (x"73",x"87",x"dd",x"fe"),
  1890 => (x"26",x"8e",x"f4",x"48"),
  1891 => (x"26",x"4c",x"26",x"4d"),
  1892 => (x"1e",x"4f",x"26",x"4b"),
  1893 => (x"86",x"f4",x"1e",x"73"),
  1894 => (x"e0",x"87",x"d1",x"fe"),
  1895 => (x"c0",x"49",x"4b",x"bf"),
  1896 => (x"02",x"99",x"c0",x"e0"),
  1897 => (x"73",x"87",x"eb",x"c0"),
  1898 => (x"9a",x"ff",x"c3",x"4a"),
  1899 => (x"97",x"cc",x"fb",x"c2"),
  1900 => (x"fb",x"c2",x"49",x"bf"),
  1901 => (x"51",x"72",x"81",x"ce"),
  1902 => (x"97",x"cc",x"fb",x"c2"),
  1903 => (x"a6",x"c4",x"48",x"bf"),
  1904 => (x"c8",x"80",x"c1",x"58"),
  1905 => (x"98",x"c7",x"58",x"a6"),
  1906 => (x"c2",x"58",x"a6",x"cc"),
  1907 => (x"c8",x"48",x"cc",x"fb"),
  1908 => (x"c8",x"fd",x"50",x"66"),
  1909 => (x"58",x"a6",x"c4",x"87"),
  1910 => (x"f4",x"87",x"c9",x"fd"),
  1911 => (x"26",x"4b",x"26",x"8e"),
  1912 => (x"fb",x"c2",x"1e",x"4f"),
  1913 => (x"cb",x"fd",x"49",x"cc"),
  1914 => (x"d3",x"f6",x"c1",x"87"),
  1915 => (x"87",x"d8",x"fc",x"49"),
  1916 => (x"26",x"87",x"e9",x"c4"),
  1917 => (x"5b",x"5e",x"0e",x"4f"),
  1918 => (x"fc",x"0e",x"5d",x"5c"),
  1919 => (x"59",x"a6",x"c4",x"86"),
  1920 => (x"c2",x"4d",x"d4",x"ff"),
  1921 => (x"fc",x"49",x"cc",x"fb"),
  1922 => (x"4b",x"70",x"87",x"f2"),
  1923 => (x"04",x"ab",x"b7",x"c0"),
  1924 => (x"c3",x"87",x"f5",x"c2"),
  1925 => (x"c9",x"05",x"ab",x"f0"),
  1926 => (x"d4",x"fb",x"c1",x"87"),
  1927 => (x"c2",x"78",x"c1",x"48"),
  1928 => (x"e0",x"c3",x"87",x"d6"),
  1929 => (x"87",x"c9",x"05",x"ab"),
  1930 => (x"48",x"d8",x"fb",x"c1"),
  1931 => (x"c7",x"c2",x"78",x"c1"),
  1932 => (x"d8",x"fb",x"c1",x"87"),
  1933 => (x"87",x"c6",x"02",x"bf"),
  1934 => (x"4c",x"a3",x"c0",x"c2"),
  1935 => (x"4c",x"73",x"87",x"c2"),
  1936 => (x"bf",x"d4",x"fb",x"c1"),
  1937 => (x"87",x"e0",x"c0",x"02"),
  1938 => (x"b7",x"c4",x"49",x"74"),
  1939 => (x"fb",x"c1",x"91",x"29"),
  1940 => (x"4a",x"74",x"81",x"dc"),
  1941 => (x"92",x"c2",x"9a",x"cf"),
  1942 => (x"30",x"72",x"48",x"c1"),
  1943 => (x"ba",x"ff",x"4a",x"70"),
  1944 => (x"98",x"69",x"48",x"72"),
  1945 => (x"87",x"db",x"79",x"70"),
  1946 => (x"b7",x"c4",x"49",x"74"),
  1947 => (x"fb",x"c1",x"91",x"29"),
  1948 => (x"4a",x"74",x"81",x"dc"),
  1949 => (x"92",x"c2",x"9a",x"cf"),
  1950 => (x"30",x"72",x"48",x"c3"),
  1951 => (x"69",x"48",x"4a",x"70"),
  1952 => (x"6e",x"79",x"70",x"b0"),
  1953 => (x"87",x"e4",x"c0",x"05"),
  1954 => (x"c8",x"48",x"d0",x"ff"),
  1955 => (x"7d",x"c5",x"78",x"e1"),
  1956 => (x"bf",x"d8",x"fb",x"c1"),
  1957 => (x"c3",x"87",x"c3",x"02"),
  1958 => (x"fb",x"c1",x"7d",x"e0"),
  1959 => (x"c3",x"02",x"bf",x"d4"),
  1960 => (x"7d",x"f0",x"c3",x"87"),
  1961 => (x"d0",x"ff",x"7d",x"73"),
  1962 => (x"78",x"e0",x"c0",x"48"),
  1963 => (x"48",x"d8",x"fb",x"c1"),
  1964 => (x"fb",x"c1",x"78",x"c0"),
  1965 => (x"78",x"c0",x"48",x"d4"),
  1966 => (x"49",x"cc",x"fb",x"c2"),
  1967 => (x"70",x"87",x"fd",x"f9"),
  1968 => (x"ab",x"b7",x"c0",x"4b"),
  1969 => (x"87",x"cb",x"fd",x"03"),
  1970 => (x"8e",x"fc",x"48",x"c0"),
  1971 => (x"4c",x"26",x"4d",x"26"),
  1972 => (x"4f",x"26",x"4b",x"26"),
  1973 => (x"00",x"00",x"00",x"00"),
  1974 => (x"00",x"00",x"00",x"00"),
  1975 => (x"00",x"00",x"00",x"00"),
  1976 => (x"34",x"34",x"34",x"34"),
  1977 => (x"34",x"34",x"34",x"34"),
  1978 => (x"34",x"34",x"34",x"34"),
  1979 => (x"34",x"34",x"34",x"34"),
  1980 => (x"34",x"34",x"34",x"34"),
  1981 => (x"34",x"34",x"34",x"34"),
  1982 => (x"34",x"34",x"34",x"34"),
  1983 => (x"34",x"34",x"34",x"34"),
  1984 => (x"34",x"34",x"34",x"34"),
  1985 => (x"34",x"34",x"34",x"34"),
  1986 => (x"34",x"34",x"34",x"34"),
  1987 => (x"34",x"34",x"34",x"34"),
  1988 => (x"34",x"34",x"34",x"34"),
  1989 => (x"34",x"34",x"34",x"34"),
  1990 => (x"34",x"34",x"34",x"34"),
  1991 => (x"72",x"4a",x"c0",x"1e"),
  1992 => (x"c1",x"91",x"c4",x"49"),
  1993 => (x"c0",x"81",x"dc",x"fb"),
  1994 => (x"d0",x"82",x"c1",x"79"),
  1995 => (x"ee",x"04",x"aa",x"b7"),
  1996 => (x"0e",x"4f",x"26",x"87"),
  1997 => (x"5d",x"5c",x"5b",x"5e"),
  1998 => (x"f7",x"4d",x"71",x"0e"),
  1999 => (x"4a",x"75",x"87",x"ee"),
  2000 => (x"92",x"2a",x"b7",x"c4"),
  2001 => (x"82",x"dc",x"fb",x"c1"),
  2002 => (x"9c",x"cf",x"4c",x"75"),
  2003 => (x"49",x"6a",x"94",x"c2"),
  2004 => (x"c3",x"2b",x"74",x"4b"),
  2005 => (x"74",x"48",x"c2",x"9b"),
  2006 => (x"ff",x"4c",x"70",x"30"),
  2007 => (x"71",x"48",x"74",x"bc"),
  2008 => (x"f6",x"7a",x"70",x"98"),
  2009 => (x"48",x"73",x"87",x"fe"),
  2010 => (x"4c",x"26",x"4d",x"26"),
  2011 => (x"4f",x"26",x"4b",x"26"),
  2012 => (x"48",x"d0",x"ff",x"1e"),
  2013 => (x"71",x"78",x"e1",x"c8"),
  2014 => (x"08",x"d4",x"ff",x"48"),
  2015 => (x"1e",x"4f",x"26",x"78"),
  2016 => (x"c8",x"48",x"d0",x"ff"),
  2017 => (x"48",x"71",x"78",x"e1"),
  2018 => (x"78",x"08",x"d4",x"ff"),
  2019 => (x"ff",x"48",x"66",x"c4"),
  2020 => (x"26",x"78",x"08",x"d4"),
  2021 => (x"4a",x"71",x"1e",x"4f"),
  2022 => (x"1e",x"49",x"66",x"c4"),
  2023 => (x"de",x"ff",x"49",x"72"),
  2024 => (x"48",x"d0",x"ff",x"87"),
  2025 => (x"fc",x"78",x"e0",x"c0"),
  2026 => (x"1e",x"4f",x"26",x"8e"),
  2027 => (x"4b",x"71",x"1e",x"73"),
  2028 => (x"1e",x"49",x"66",x"c8"),
  2029 => (x"e0",x"c1",x"4a",x"73"),
  2030 => (x"d8",x"ff",x"49",x"a2"),
  2031 => (x"26",x"8e",x"fc",x"87"),
  2032 => (x"1e",x"4f",x"26",x"4b"),
  2033 => (x"c8",x"48",x"d0",x"ff"),
  2034 => (x"48",x"71",x"78",x"c9"),
  2035 => (x"78",x"08",x"d4",x"ff"),
  2036 => (x"71",x"1e",x"4f",x"26"),
  2037 => (x"87",x"eb",x"49",x"4a"),
  2038 => (x"c8",x"48",x"d0",x"ff"),
  2039 => (x"1e",x"4f",x"26",x"78"),
  2040 => (x"4b",x"71",x"1e",x"73"),
  2041 => (x"bf",x"e4",x"fb",x"c2"),
  2042 => (x"c2",x"87",x"c3",x"02"),
  2043 => (x"d0",x"ff",x"87",x"eb"),
  2044 => (x"78",x"c9",x"c8",x"48"),
  2045 => (x"e0",x"c0",x"48",x"73"),
  2046 => (x"08",x"d4",x"ff",x"b0"),
  2047 => (x"d8",x"fb",x"c2",x"78"),
  2048 => (x"c8",x"78",x"c0",x"48"),
  2049 => (x"87",x"c5",x"02",x"66"),
  2050 => (x"c2",x"49",x"ff",x"c3"),
  2051 => (x"c2",x"49",x"c0",x"87"),
  2052 => (x"cc",x"59",x"e0",x"fb"),
  2053 => (x"87",x"c6",x"02",x"66"),
  2054 => (x"4a",x"d5",x"d5",x"c5"),
  2055 => (x"ff",x"cf",x"87",x"c4"),
  2056 => (x"fb",x"c2",x"4a",x"ff"),
  2057 => (x"fb",x"c2",x"5a",x"e4"),
  2058 => (x"78",x"c1",x"48",x"e4"),
  2059 => (x"4f",x"26",x"4b",x"26"),
  2060 => (x"5c",x"5b",x"5e",x"0e"),
  2061 => (x"4d",x"71",x"0e",x"5d"),
  2062 => (x"bf",x"e0",x"fb",x"c2"),
  2063 => (x"02",x"9d",x"75",x"4b"),
  2064 => (x"c8",x"49",x"87",x"cb"),
  2065 => (x"d8",x"ff",x"c1",x"91"),
  2066 => (x"c4",x"82",x"71",x"4a"),
  2067 => (x"d8",x"c3",x"c2",x"87"),
  2068 => (x"12",x"4c",x"c0",x"4a"),
  2069 => (x"c2",x"99",x"73",x"49"),
  2070 => (x"48",x"bf",x"dc",x"fb"),
  2071 => (x"d4",x"ff",x"b8",x"71"),
  2072 => (x"b7",x"c1",x"78",x"08"),
  2073 => (x"b7",x"c8",x"84",x"2b"),
  2074 => (x"87",x"e7",x"04",x"ac"),
  2075 => (x"bf",x"d8",x"fb",x"c2"),
  2076 => (x"c2",x"80",x"c8",x"48"),
  2077 => (x"26",x"58",x"dc",x"fb"),
  2078 => (x"26",x"4c",x"26",x"4d"),
  2079 => (x"1e",x"4f",x"26",x"4b"),
  2080 => (x"4b",x"71",x"1e",x"73"),
  2081 => (x"02",x"9a",x"4a",x"13"),
  2082 => (x"49",x"72",x"87",x"cb"),
  2083 => (x"13",x"87",x"e1",x"fe"),
  2084 => (x"f5",x"05",x"9a",x"4a"),
  2085 => (x"26",x"4b",x"26",x"87"),
  2086 => (x"fb",x"c2",x"1e",x"4f"),
  2087 => (x"c2",x"49",x"bf",x"d8"),
  2088 => (x"c1",x"48",x"d8",x"fb"),
  2089 => (x"c0",x"c4",x"78",x"a1"),
  2090 => (x"db",x"03",x"a9",x"b7"),
  2091 => (x"48",x"d4",x"ff",x"87"),
  2092 => (x"bf",x"dc",x"fb",x"c2"),
  2093 => (x"d8",x"fb",x"c2",x"78"),
  2094 => (x"fb",x"c2",x"49",x"bf"),
  2095 => (x"a1",x"c1",x"48",x"d8"),
  2096 => (x"b7",x"c0",x"c4",x"78"),
  2097 => (x"87",x"e5",x"04",x"a9"),
  2098 => (x"c8",x"48",x"d0",x"ff"),
  2099 => (x"e4",x"fb",x"c2",x"78"),
  2100 => (x"26",x"78",x"c0",x"48"),
  2101 => (x"00",x"00",x"00",x"4f"),
  2102 => (x"00",x"00",x"00",x"00"),
  2103 => (x"00",x"00",x"00",x"00"),
  2104 => (x"5f",x"00",x"00",x"00"),
  2105 => (x"00",x"00",x"00",x"5f"),
  2106 => (x"00",x"03",x"03",x"00"),
  2107 => (x"00",x"00",x"03",x"03"),
  2108 => (x"14",x"7f",x"7f",x"14"),
  2109 => (x"00",x"14",x"7f",x"7f"),
  2110 => (x"6b",x"2e",x"24",x"00"),
  2111 => (x"00",x"12",x"3a",x"6b"),
  2112 => (x"18",x"36",x"6a",x"4c"),
  2113 => (x"00",x"32",x"56",x"6c"),
  2114 => (x"59",x"4f",x"7e",x"30"),
  2115 => (x"40",x"68",x"3a",x"77"),
  2116 => (x"07",x"04",x"00",x"00"),
  2117 => (x"00",x"00",x"00",x"03"),
  2118 => (x"3e",x"1c",x"00",x"00"),
  2119 => (x"00",x"00",x"41",x"63"),
  2120 => (x"63",x"41",x"00",x"00"),
  2121 => (x"00",x"00",x"1c",x"3e"),
  2122 => (x"1c",x"3e",x"2a",x"08"),
  2123 => (x"08",x"2a",x"3e",x"1c"),
  2124 => (x"3e",x"08",x"08",x"00"),
  2125 => (x"00",x"08",x"08",x"3e"),
  2126 => (x"e0",x"80",x"00",x"00"),
  2127 => (x"00",x"00",x"00",x"60"),
  2128 => (x"08",x"08",x"08",x"00"),
  2129 => (x"00",x"08",x"08",x"08"),
  2130 => (x"60",x"00",x"00",x"00"),
  2131 => (x"00",x"00",x"00",x"60"),
  2132 => (x"18",x"30",x"60",x"40"),
  2133 => (x"01",x"03",x"06",x"0c"),
  2134 => (x"59",x"7f",x"3e",x"00"),
  2135 => (x"00",x"3e",x"7f",x"4d"),
  2136 => (x"7f",x"06",x"04",x"00"),
  2137 => (x"00",x"00",x"00",x"7f"),
  2138 => (x"71",x"63",x"42",x"00"),
  2139 => (x"00",x"46",x"4f",x"59"),
  2140 => (x"49",x"63",x"22",x"00"),
  2141 => (x"00",x"36",x"7f",x"49"),
  2142 => (x"13",x"16",x"1c",x"18"),
  2143 => (x"00",x"10",x"7f",x"7f"),
  2144 => (x"45",x"67",x"27",x"00"),
  2145 => (x"00",x"39",x"7d",x"45"),
  2146 => (x"4b",x"7e",x"3c",x"00"),
  2147 => (x"00",x"30",x"79",x"49"),
  2148 => (x"71",x"01",x"01",x"00"),
  2149 => (x"00",x"07",x"0f",x"79"),
  2150 => (x"49",x"7f",x"36",x"00"),
  2151 => (x"00",x"36",x"7f",x"49"),
  2152 => (x"49",x"4f",x"06",x"00"),
  2153 => (x"00",x"1e",x"3f",x"69"),
  2154 => (x"66",x"00",x"00",x"00"),
  2155 => (x"00",x"00",x"00",x"66"),
  2156 => (x"e6",x"80",x"00",x"00"),
  2157 => (x"00",x"00",x"00",x"66"),
  2158 => (x"14",x"08",x"08",x"00"),
  2159 => (x"00",x"22",x"22",x"14"),
  2160 => (x"14",x"14",x"14",x"00"),
  2161 => (x"00",x"14",x"14",x"14"),
  2162 => (x"14",x"22",x"22",x"00"),
  2163 => (x"00",x"08",x"08",x"14"),
  2164 => (x"51",x"03",x"02",x"00"),
  2165 => (x"00",x"06",x"0f",x"59"),
  2166 => (x"5d",x"41",x"7f",x"3e"),
  2167 => (x"00",x"1e",x"1f",x"55"),
  2168 => (x"09",x"7f",x"7e",x"00"),
  2169 => (x"00",x"7e",x"7f",x"09"),
  2170 => (x"49",x"7f",x"7f",x"00"),
  2171 => (x"00",x"36",x"7f",x"49"),
  2172 => (x"63",x"3e",x"1c",x"00"),
  2173 => (x"00",x"41",x"41",x"41"),
  2174 => (x"41",x"7f",x"7f",x"00"),
  2175 => (x"00",x"1c",x"3e",x"63"),
  2176 => (x"49",x"7f",x"7f",x"00"),
  2177 => (x"00",x"41",x"41",x"49"),
  2178 => (x"09",x"7f",x"7f",x"00"),
  2179 => (x"00",x"01",x"01",x"09"),
  2180 => (x"41",x"7f",x"3e",x"00"),
  2181 => (x"00",x"7a",x"7b",x"49"),
  2182 => (x"08",x"7f",x"7f",x"00"),
  2183 => (x"00",x"7f",x"7f",x"08"),
  2184 => (x"7f",x"41",x"00",x"00"),
  2185 => (x"00",x"00",x"41",x"7f"),
  2186 => (x"40",x"60",x"20",x"00"),
  2187 => (x"00",x"3f",x"7f",x"40"),
  2188 => (x"1c",x"08",x"7f",x"7f"),
  2189 => (x"00",x"41",x"63",x"36"),
  2190 => (x"40",x"7f",x"7f",x"00"),
  2191 => (x"00",x"40",x"40",x"40"),
  2192 => (x"0c",x"06",x"7f",x"7f"),
  2193 => (x"00",x"7f",x"7f",x"06"),
  2194 => (x"0c",x"06",x"7f",x"7f"),
  2195 => (x"00",x"7f",x"7f",x"18"),
  2196 => (x"41",x"7f",x"3e",x"00"),
  2197 => (x"00",x"3e",x"7f",x"41"),
  2198 => (x"09",x"7f",x"7f",x"00"),
  2199 => (x"00",x"06",x"0f",x"09"),
  2200 => (x"61",x"41",x"7f",x"3e"),
  2201 => (x"00",x"40",x"7e",x"7f"),
  2202 => (x"09",x"7f",x"7f",x"00"),
  2203 => (x"00",x"66",x"7f",x"19"),
  2204 => (x"4d",x"6f",x"26",x"00"),
  2205 => (x"00",x"32",x"7b",x"59"),
  2206 => (x"7f",x"01",x"01",x"00"),
  2207 => (x"00",x"01",x"01",x"7f"),
  2208 => (x"40",x"7f",x"3f",x"00"),
  2209 => (x"00",x"3f",x"7f",x"40"),
  2210 => (x"70",x"3f",x"0f",x"00"),
  2211 => (x"00",x"0f",x"3f",x"70"),
  2212 => (x"18",x"30",x"7f",x"7f"),
  2213 => (x"00",x"7f",x"7f",x"30"),
  2214 => (x"1c",x"36",x"63",x"41"),
  2215 => (x"41",x"63",x"36",x"1c"),
  2216 => (x"7c",x"06",x"03",x"01"),
  2217 => (x"01",x"03",x"06",x"7c"),
  2218 => (x"4d",x"59",x"71",x"61"),
  2219 => (x"00",x"41",x"43",x"47"),
  2220 => (x"7f",x"7f",x"00",x"00"),
  2221 => (x"00",x"00",x"41",x"41"),
  2222 => (x"0c",x"06",x"03",x"01"),
  2223 => (x"40",x"60",x"30",x"18"),
  2224 => (x"41",x"41",x"00",x"00"),
  2225 => (x"00",x"00",x"7f",x"7f"),
  2226 => (x"03",x"06",x"0c",x"08"),
  2227 => (x"00",x"08",x"0c",x"06"),
  2228 => (x"80",x"80",x"80",x"80"),
  2229 => (x"00",x"80",x"80",x"80"),
  2230 => (x"03",x"00",x"00",x"00"),
  2231 => (x"00",x"00",x"04",x"07"),
  2232 => (x"54",x"74",x"20",x"00"),
  2233 => (x"00",x"78",x"7c",x"54"),
  2234 => (x"44",x"7f",x"7f",x"00"),
  2235 => (x"00",x"38",x"7c",x"44"),
  2236 => (x"44",x"7c",x"38",x"00"),
  2237 => (x"00",x"00",x"44",x"44"),
  2238 => (x"44",x"7c",x"38",x"00"),
  2239 => (x"00",x"7f",x"7f",x"44"),
  2240 => (x"54",x"7c",x"38",x"00"),
  2241 => (x"00",x"18",x"5c",x"54"),
  2242 => (x"7f",x"7e",x"04",x"00"),
  2243 => (x"00",x"00",x"05",x"05"),
  2244 => (x"a4",x"bc",x"18",x"00"),
  2245 => (x"00",x"7c",x"fc",x"a4"),
  2246 => (x"04",x"7f",x"7f",x"00"),
  2247 => (x"00",x"78",x"7c",x"04"),
  2248 => (x"3d",x"00",x"00",x"00"),
  2249 => (x"00",x"00",x"40",x"7d"),
  2250 => (x"80",x"80",x"80",x"00"),
  2251 => (x"00",x"00",x"7d",x"fd"),
  2252 => (x"10",x"7f",x"7f",x"00"),
  2253 => (x"00",x"44",x"6c",x"38"),
  2254 => (x"3f",x"00",x"00",x"00"),
  2255 => (x"00",x"00",x"40",x"7f"),
  2256 => (x"18",x"0c",x"7c",x"7c"),
  2257 => (x"00",x"78",x"7c",x"0c"),
  2258 => (x"04",x"7c",x"7c",x"00"),
  2259 => (x"00",x"78",x"7c",x"04"),
  2260 => (x"44",x"7c",x"38",x"00"),
  2261 => (x"00",x"38",x"7c",x"44"),
  2262 => (x"24",x"fc",x"fc",x"00"),
  2263 => (x"00",x"18",x"3c",x"24"),
  2264 => (x"24",x"3c",x"18",x"00"),
  2265 => (x"00",x"fc",x"fc",x"24"),
  2266 => (x"04",x"7c",x"7c",x"00"),
  2267 => (x"00",x"08",x"0c",x"04"),
  2268 => (x"54",x"5c",x"48",x"00"),
  2269 => (x"00",x"20",x"74",x"54"),
  2270 => (x"7f",x"3f",x"04",x"00"),
  2271 => (x"00",x"00",x"44",x"44"),
  2272 => (x"40",x"7c",x"3c",x"00"),
  2273 => (x"00",x"7c",x"7c",x"40"),
  2274 => (x"60",x"3c",x"1c",x"00"),
  2275 => (x"00",x"1c",x"3c",x"60"),
  2276 => (x"30",x"60",x"7c",x"3c"),
  2277 => (x"00",x"3c",x"7c",x"60"),
  2278 => (x"10",x"38",x"6c",x"44"),
  2279 => (x"00",x"44",x"6c",x"38"),
  2280 => (x"e0",x"bc",x"1c",x"00"),
  2281 => (x"00",x"1c",x"3c",x"60"),
  2282 => (x"74",x"64",x"44",x"00"),
  2283 => (x"00",x"44",x"4c",x"5c"),
  2284 => (x"3e",x"08",x"08",x"00"),
  2285 => (x"00",x"41",x"41",x"77"),
  2286 => (x"7f",x"00",x"00",x"00"),
  2287 => (x"00",x"00",x"00",x"7f"),
  2288 => (x"77",x"41",x"41",x"00"),
  2289 => (x"00",x"08",x"08",x"3e"),
  2290 => (x"03",x"01",x"01",x"02"),
  2291 => (x"00",x"01",x"02",x"02"),
  2292 => (x"7f",x"7f",x"7f",x"7f"),
  2293 => (x"00",x"7f",x"7f",x"7f"),
  2294 => (x"1c",x"1c",x"08",x"08"),
  2295 => (x"7f",x"7f",x"3e",x"3e"),
  2296 => (x"3e",x"3e",x"7f",x"7f"),
  2297 => (x"08",x"08",x"1c",x"1c"),
  2298 => (x"7c",x"18",x"10",x"00"),
  2299 => (x"00",x"10",x"18",x"7c"),
  2300 => (x"7c",x"30",x"10",x"00"),
  2301 => (x"00",x"10",x"30",x"7c"),
  2302 => (x"60",x"60",x"30",x"10"),
  2303 => (x"00",x"06",x"1e",x"78"),
  2304 => (x"18",x"3c",x"66",x"42"),
  2305 => (x"00",x"42",x"66",x"3c"),
  2306 => (x"c2",x"6a",x"38",x"78"),
  2307 => (x"00",x"38",x"6c",x"c6"),
  2308 => (x"60",x"00",x"00",x"60"),
  2309 => (x"00",x"60",x"00",x"00"),
  2310 => (x"5c",x"5b",x"5e",x"0e"),
  2311 => (x"86",x"fc",x"0e",x"5d"),
  2312 => (x"c2",x"59",x"a6",x"c4"),
  2313 => (x"4c",x"bf",x"ec",x"fb"),
  2314 => (x"1e",x"c0",x"4b",x"c0"),
  2315 => (x"02",x"ab",x"66",x"c4"),
  2316 => (x"4d",x"c0",x"87",x"c4"),
  2317 => (x"4d",x"c1",x"87",x"c2"),
  2318 => (x"49",x"73",x"1e",x"75"),
  2319 => (x"c8",x"87",x"e0",x"ee"),
  2320 => (x"49",x"e0",x"c0",x"86"),
  2321 => (x"c4",x"87",x"e9",x"ef"),
  2322 => (x"49",x"6a",x"4a",x"a4"),
  2323 => (x"f1",x"87",x"f0",x"f0"),
  2324 => (x"84",x"cc",x"87",x"c7"),
  2325 => (x"b7",x"c8",x"83",x"c1"),
  2326 => (x"cd",x"ff",x"04",x"ab"),
  2327 => (x"26",x"8e",x"fc",x"87"),
  2328 => (x"26",x"4c",x"26",x"4d"),
  2329 => (x"1e",x"4f",x"26",x"4b"),
  2330 => (x"fb",x"c2",x"4a",x"71"),
  2331 => (x"fb",x"c2",x"5a",x"f0"),
  2332 => (x"78",x"c7",x"48",x"f0"),
  2333 => (x"87",x"e0",x"fe",x"49"),
  2334 => (x"73",x"1e",x"4f",x"26"),
  2335 => (x"fc",x"4b",x"71",x"1e"),
  2336 => (x"73",x"0b",x"7b",x"0b"),
  2337 => (x"c1",x"9a",x"c1",x"4a"),
  2338 => (x"ed",x"49",x"a2",x"c0"),
  2339 => (x"df",x"c2",x"87",x"c4"),
  2340 => (x"4b",x"26",x"5b",x"f0"),
  2341 => (x"71",x"1e",x"4f",x"26"),
  2342 => (x"1e",x"66",x"c4",x"4a"),
  2343 => (x"ca",x"ec",x"49",x"72"),
  2344 => (x"26",x"8e",x"fc",x"87"),
  2345 => (x"d4",x"ff",x"1e",x"4f"),
  2346 => (x"78",x"ff",x"c3",x"48"),
  2347 => (x"c0",x"48",x"d0",x"ff"),
  2348 => (x"d4",x"ff",x"78",x"e1"),
  2349 => (x"71",x"78",x"c1",x"48"),
  2350 => (x"ff",x"30",x"c4",x"48"),
  2351 => (x"ff",x"78",x"08",x"d4"),
  2352 => (x"e0",x"c0",x"48",x"d0"),
  2353 => (x"0e",x"4f",x"26",x"78"),
  2354 => (x"5d",x"5c",x"5b",x"5e"),
  2355 => (x"c8",x"86",x"ec",x"0e"),
  2356 => (x"78",x"c0",x"48",x"a6"),
  2357 => (x"bf",x"ec",x"80",x"c4"),
  2358 => (x"c2",x"80",x"f8",x"78"),
  2359 => (x"78",x"bf",x"ec",x"fb"),
  2360 => (x"bf",x"f4",x"fb",x"c2"),
  2361 => (x"4d",x"bf",x"e8",x"4c"),
  2362 => (x"bf",x"ec",x"df",x"c2"),
  2363 => (x"87",x"c5",x"e4",x"49"),
  2364 => (x"fe",x"e8",x"49",x"c7"),
  2365 => (x"c2",x"49",x"70",x"87"),
  2366 => (x"87",x"d0",x"05",x"99"),
  2367 => (x"bf",x"e4",x"df",x"c2"),
  2368 => (x"cc",x"b9",x"ff",x"49"),
  2369 => (x"99",x"c1",x"99",x"66"),
  2370 => (x"87",x"cd",x"c2",x"02"),
  2371 => (x"ff",x"48",x"a6",x"c8"),
  2372 => (x"c7",x"78",x"bf",x"c8"),
  2373 => (x"87",x"db",x"e8",x"49"),
  2374 => (x"a6",x"c4",x"49",x"70"),
  2375 => (x"05",x"99",x"71",x"5c"),
  2376 => (x"66",x"cc",x"87",x"ce"),
  2377 => (x"c4",x"99",x"c1",x"49"),
  2378 => (x"99",x"71",x"5c",x"a6"),
  2379 => (x"87",x"c4",x"c1",x"02"),
  2380 => (x"c8",x"4c",x"c8",x"ff"),
  2381 => (x"a6",x"cc",x"4b",x"66"),
  2382 => (x"78",x"bf",x"ec",x"48"),
  2383 => (x"cc",x"87",x"f6",x"e2"),
  2384 => (x"48",x"6c",x"5b",x"a6"),
  2385 => (x"a6",x"d4",x"88",x"73"),
  2386 => (x"a8",x"e8",x"cf",x"58"),
  2387 => (x"c2",x"87",x"d1",x"06"),
  2388 => (x"49",x"bf",x"e0",x"df"),
  2389 => (x"df",x"c2",x"b9",x"c1"),
  2390 => (x"fd",x"71",x"59",x"e4"),
  2391 => (x"4b",x"6c",x"87",x"c7"),
  2392 => (x"ce",x"e7",x"49",x"c7"),
  2393 => (x"05",x"98",x"70",x"87"),
  2394 => (x"cc",x"87",x"cb",x"ff"),
  2395 => (x"99",x"c1",x"49",x"66"),
  2396 => (x"87",x"c2",x"ff",x"05"),
  2397 => (x"df",x"c2",x"4c",x"6e"),
  2398 => (x"c1",x"4a",x"bf",x"ec"),
  2399 => (x"f0",x"df",x"c2",x"ba"),
  2400 => (x"7a",x"0a",x"fc",x"5a"),
  2401 => (x"c1",x"9a",x"c1",x"0a"),
  2402 => (x"e9",x"49",x"a2",x"c0"),
  2403 => (x"da",x"c1",x"87",x"c4"),
  2404 => (x"87",x"df",x"e6",x"49"),
  2405 => (x"c1",x"48",x"a6",x"c8"),
  2406 => (x"e4",x"df",x"c2",x"78"),
  2407 => (x"78",x"66",x"cc",x"48"),
  2408 => (x"bf",x"ec",x"df",x"c2"),
  2409 => (x"87",x"c7",x"c1",x"05"),
  2410 => (x"4b",x"c0",x"c0",x"c8"),
  2411 => (x"7e",x"d0",x"df",x"c2"),
  2412 => (x"49",x"14",x"4c",x"6e"),
  2413 => (x"70",x"87",x"fc",x"e5"),
  2414 => (x"c2",x"c0",x"02",x"98"),
  2415 => (x"c1",x"b5",x"73",x"87"),
  2416 => (x"ff",x"05",x"2b",x"b7"),
  2417 => (x"49",x"75",x"87",x"ec"),
  2418 => (x"71",x"99",x"ff",x"c3"),
  2419 => (x"fb",x"49",x"c0",x"1e"),
  2420 => (x"49",x"75",x"87",x"c4"),
  2421 => (x"71",x"29",x"b7",x"c8"),
  2422 => (x"fa",x"49",x"c1",x"1e"),
  2423 => (x"86",x"c8",x"87",x"f8"),
  2424 => (x"e5",x"49",x"fd",x"c3"),
  2425 => (x"fa",x"c3",x"87",x"cd"),
  2426 => (x"87",x"c7",x"e5",x"49"),
  2427 => (x"75",x"87",x"d2",x"c7"),
  2428 => (x"99",x"ff",x"c3",x"49"),
  2429 => (x"71",x"2d",x"b7",x"c8"),
  2430 => (x"02",x"9d",x"75",x"b5"),
  2431 => (x"ff",x"87",x"e0",x"c0"),
  2432 => (x"6e",x"7e",x"bf",x"c8"),
  2433 => (x"e8",x"df",x"c2",x"49"),
  2434 => (x"e0",x"c2",x"89",x"bf"),
  2435 => (x"c5",x"c0",x"03",x"a9"),
  2436 => (x"c0",x"4d",x"c0",x"87"),
  2437 => (x"df",x"c2",x"87",x"cf"),
  2438 => (x"78",x"6e",x"48",x"e8"),
  2439 => (x"c2",x"87",x"c6",x"c0"),
  2440 => (x"c0",x"48",x"e8",x"df"),
  2441 => (x"c8",x"49",x"75",x"78"),
  2442 => (x"ce",x"c0",x"05",x"99"),
  2443 => (x"49",x"f5",x"c3",x"87"),
  2444 => (x"70",x"87",x"c0",x"e4"),
  2445 => (x"02",x"99",x"c2",x"49"),
  2446 => (x"c2",x"87",x"eb",x"c0"),
  2447 => (x"02",x"bf",x"f0",x"fb"),
  2448 => (x"48",x"87",x"ca",x"c0"),
  2449 => (x"fb",x"c2",x"88",x"c1"),
  2450 => (x"d4",x"c0",x"58",x"f4"),
  2451 => (x"48",x"66",x"c4",x"87"),
  2452 => (x"c4",x"80",x"e0",x"c1"),
  2453 => (x"bf",x"6e",x"58",x"a6"),
  2454 => (x"87",x"c5",x"c0",x"02"),
  2455 => (x"73",x"49",x"ff",x"4b"),
  2456 => (x"48",x"a6",x"c8",x"0f"),
  2457 => (x"49",x"75",x"78",x"c1"),
  2458 => (x"c0",x"05",x"99",x"c4"),
  2459 => (x"f2",x"c3",x"87",x"ce"),
  2460 => (x"87",x"ff",x"e2",x"49"),
  2461 => (x"99",x"c2",x"49",x"70"),
  2462 => (x"87",x"f2",x"c0",x"02"),
  2463 => (x"bf",x"f0",x"fb",x"c2"),
  2464 => (x"c7",x"48",x"6e",x"7e"),
  2465 => (x"c0",x"03",x"a8",x"b7"),
  2466 => (x"48",x"6e",x"87",x"cb"),
  2467 => (x"fb",x"c2",x"80",x"c1"),
  2468 => (x"d4",x"c0",x"58",x"f4"),
  2469 => (x"48",x"66",x"c4",x"87"),
  2470 => (x"c4",x"80",x"e0",x"c1"),
  2471 => (x"bf",x"6e",x"58",x"a6"),
  2472 => (x"87",x"c5",x"c0",x"02"),
  2473 => (x"73",x"49",x"fe",x"4b"),
  2474 => (x"48",x"a6",x"c8",x"0f"),
  2475 => (x"fd",x"c3",x"78",x"c1"),
  2476 => (x"87",x"ff",x"e1",x"49"),
  2477 => (x"99",x"c2",x"49",x"70"),
  2478 => (x"87",x"e6",x"c0",x"02"),
  2479 => (x"bf",x"f0",x"fb",x"c2"),
  2480 => (x"87",x"c9",x"c0",x"02"),
  2481 => (x"48",x"f0",x"fb",x"c2"),
  2482 => (x"d0",x"c0",x"78",x"c0"),
  2483 => (x"4a",x"66",x"c4",x"87"),
  2484 => (x"6a",x"82",x"e0",x"c1"),
  2485 => (x"87",x"c5",x"c0",x"02"),
  2486 => (x"73",x"49",x"fd",x"4b"),
  2487 => (x"48",x"a6",x"c8",x"0f"),
  2488 => (x"fa",x"c3",x"78",x"c1"),
  2489 => (x"87",x"cb",x"e1",x"49"),
  2490 => (x"99",x"c2",x"49",x"70"),
  2491 => (x"87",x"ee",x"c0",x"02"),
  2492 => (x"bf",x"f0",x"fb",x"c2"),
  2493 => (x"a8",x"b7",x"c7",x"48"),
  2494 => (x"87",x"c9",x"c0",x"03"),
  2495 => (x"48",x"f0",x"fb",x"c2"),
  2496 => (x"d4",x"c0",x"78",x"c7"),
  2497 => (x"48",x"66",x"c4",x"87"),
  2498 => (x"c4",x"80",x"e0",x"c1"),
  2499 => (x"bf",x"6e",x"58",x"a6"),
  2500 => (x"87",x"c5",x"c0",x"02"),
  2501 => (x"73",x"49",x"fc",x"4b"),
  2502 => (x"48",x"a6",x"c8",x"0f"),
  2503 => (x"48",x"75",x"78",x"c1"),
  2504 => (x"c4",x"98",x"f0",x"c3"),
  2505 => (x"98",x"70",x"58",x"a6"),
  2506 => (x"87",x"ce",x"c0",x"05"),
  2507 => (x"e0",x"49",x"da",x"c1"),
  2508 => (x"49",x"70",x"87",x"c1"),
  2509 => (x"c1",x"02",x"99",x"c2"),
  2510 => (x"05",x"6e",x"87",x"ca"),
  2511 => (x"c1",x"87",x"cd",x"c0"),
  2512 => (x"df",x"ff",x"49",x"da"),
  2513 => (x"98",x"70",x"87",x"ed"),
  2514 => (x"87",x"e8",x"c0",x"02"),
  2515 => (x"4b",x"49",x"bf",x"e8"),
  2516 => (x"c8",x"9b",x"ff",x"c3"),
  2517 => (x"b3",x"71",x"29",x"b7"),
  2518 => (x"87",x"d9",x"da",x"ff"),
  2519 => (x"f0",x"c3",x"49",x"73"),
  2520 => (x"05",x"99",x"71",x"99"),
  2521 => (x"c1",x"87",x"e5",x"ff"),
  2522 => (x"df",x"ff",x"49",x"da"),
  2523 => (x"98",x"70",x"87",x"c5"),
  2524 => (x"87",x"d8",x"ff",x"05"),
  2525 => (x"bf",x"f0",x"fb",x"c2"),
  2526 => (x"93",x"cc",x"4b",x"49"),
  2527 => (x"6b",x"83",x"66",x"c4"),
  2528 => (x"0f",x"73",x"71",x"4b"),
  2529 => (x"c0",x"02",x"9c",x"74"),
  2530 => (x"02",x"6c",x"87",x"e9"),
  2531 => (x"6c",x"87",x"e4",x"c0"),
  2532 => (x"de",x"de",x"ff",x"49"),
  2533 => (x"c1",x"49",x"70",x"87"),
  2534 => (x"cb",x"c0",x"02",x"99"),
  2535 => (x"4b",x"a4",x"c4",x"87"),
  2536 => (x"bf",x"f0",x"fb",x"c2"),
  2537 => (x"0f",x"4b",x"6b",x"49"),
  2538 => (x"c0",x"02",x"84",x"c8"),
  2539 => (x"05",x"6c",x"87",x"c5"),
  2540 => (x"c8",x"87",x"dc",x"ff"),
  2541 => (x"c8",x"c0",x"02",x"66"),
  2542 => (x"f0",x"fb",x"c2",x"87"),
  2543 => (x"d7",x"f1",x"49",x"bf"),
  2544 => (x"26",x"8e",x"ec",x"87"),
  2545 => (x"26",x"4c",x"26",x"4d"),
  2546 => (x"00",x"4f",x"26",x"4b"),
  2547 => (x"00",x"00",x"00",x"10"),
  2548 => (x"14",x"11",x"12",x"58"),
  2549 => (x"23",x"1c",x"1b",x"1d"),
  2550 => (x"94",x"91",x"59",x"5a"),
  2551 => (x"f4",x"eb",x"f2",x"f5"),
  2552 => (x"00",x"00",x"00",x"00"),
  2553 => (x"00",x"00",x"00",x"00"),
  2554 => (x"00",x"00",x"00",x"00"),
  2555 => (x"00",x"00",x"00",x"00"),
  2556 => (x"5c",x"5b",x"5e",x"0e"),
  2557 => (x"4b",x"71",x"0e",x"5d"),
  2558 => (x"d0",x"4c",x"d4",x"ff"),
  2559 => (x"78",x"c0",x"48",x"66"),
  2560 => (x"dd",x"ff",x"49",x"d6"),
  2561 => (x"ff",x"c3",x"87",x"ea"),
  2562 => (x"c3",x"49",x"6c",x"7c"),
  2563 => (x"4d",x"71",x"99",x"ff"),
  2564 => (x"99",x"f0",x"c3",x"49"),
  2565 => (x"05",x"a9",x"e0",x"c1"),
  2566 => (x"ff",x"c3",x"87",x"cb"),
  2567 => (x"c3",x"48",x"6c",x"7c"),
  2568 => (x"08",x"66",x"d0",x"98"),
  2569 => (x"7c",x"ff",x"c3",x"78"),
  2570 => (x"c8",x"49",x"4a",x"6c"),
  2571 => (x"7c",x"ff",x"c3",x"31"),
  2572 => (x"b2",x"71",x"4a",x"6c"),
  2573 => (x"31",x"c8",x"49",x"72"),
  2574 => (x"6c",x"7c",x"ff",x"c3"),
  2575 => (x"72",x"b2",x"71",x"4a"),
  2576 => (x"c3",x"31",x"c8",x"49"),
  2577 => (x"4a",x"6c",x"7c",x"ff"),
  2578 => (x"d0",x"ff",x"b2",x"71"),
  2579 => (x"78",x"e0",x"c0",x"48"),
  2580 => (x"c2",x"02",x"9b",x"73"),
  2581 => (x"75",x"7b",x"72",x"87"),
  2582 => (x"26",x"4d",x"26",x"48"),
  2583 => (x"26",x"4b",x"26",x"4c"),
  2584 => (x"4f",x"26",x"1e",x"4f"),
  2585 => (x"5c",x"5b",x"5e",x"0e"),
  2586 => (x"76",x"86",x"f8",x"0e"),
  2587 => (x"80",x"c4",x"48",x"1e"),
  2588 => (x"fb",x"fd",x"49",x"70"),
  2589 => (x"70",x"86",x"c4",x"87"),
  2590 => (x"c3",x"48",x"6e",x"4b"),
  2591 => (x"f4",x"c2",x"01",x"a8"),
  2592 => (x"c3",x"4a",x"73",x"87"),
  2593 => (x"d0",x"c1",x"9a",x"f0"),
  2594 => (x"87",x"c7",x"02",x"aa"),
  2595 => (x"05",x"aa",x"e0",x"c1"),
  2596 => (x"73",x"87",x"e2",x"c2"),
  2597 => (x"02",x"99",x"c8",x"49"),
  2598 => (x"c4",x"ff",x"87",x"c3"),
  2599 => (x"c3",x"4c",x"73",x"87"),
  2600 => (x"05",x"ac",x"c2",x"9c"),
  2601 => (x"c4",x"87",x"c4",x"c1"),
  2602 => (x"31",x"c9",x"49",x"66"),
  2603 => (x"66",x"c4",x"1e",x"71"),
  2604 => (x"92",x"cc",x"c1",x"4a"),
  2605 => (x"49",x"f8",x"fb",x"c2"),
  2606 => (x"cc",x"fe",x"81",x"72"),
  2607 => (x"49",x"d8",x"87",x"fe"),
  2608 => (x"87",x"ec",x"da",x"ff"),
  2609 => (x"c2",x"1e",x"c0",x"c8"),
  2610 => (x"fd",x"49",x"f0",x"e8"),
  2611 => (x"ff",x"87",x"d0",x"e6"),
  2612 => (x"e0",x"c0",x"48",x"d0"),
  2613 => (x"f0",x"e8",x"c2",x"78"),
  2614 => (x"4a",x"66",x"cc",x"1e"),
  2615 => (x"c2",x"92",x"cc",x"c1"),
  2616 => (x"72",x"49",x"f8",x"fb"),
  2617 => (x"d4",x"cb",x"fe",x"81"),
  2618 => (x"c1",x"86",x"cc",x"87"),
  2619 => (x"c4",x"c1",x"05",x"ac"),
  2620 => (x"49",x"66",x"c4",x"87"),
  2621 => (x"1e",x"71",x"31",x"c9"),
  2622 => (x"c1",x"4a",x"66",x"c4"),
  2623 => (x"fb",x"c2",x"92",x"cc"),
  2624 => (x"81",x"72",x"49",x"f8"),
  2625 => (x"87",x"f4",x"cb",x"fe"),
  2626 => (x"1e",x"f0",x"e8",x"c2"),
  2627 => (x"c1",x"4a",x"66",x"c8"),
  2628 => (x"fb",x"c2",x"92",x"cc"),
  2629 => (x"81",x"72",x"49",x"f8"),
  2630 => (x"87",x"e2",x"c9",x"fe"),
  2631 => (x"d9",x"ff",x"49",x"d7"),
  2632 => (x"c0",x"c8",x"87",x"ce"),
  2633 => (x"f0",x"e8",x"c2",x"1e"),
  2634 => (x"cf",x"e4",x"fd",x"49"),
  2635 => (x"ff",x"86",x"cc",x"87"),
  2636 => (x"e0",x"c0",x"48",x"d0"),
  2637 => (x"26",x"8e",x"f8",x"78"),
  2638 => (x"26",x"4b",x"26",x"4c"),
  2639 => (x"4a",x"71",x"1e",x"4f"),
  2640 => (x"03",x"aa",x"b7",x"c4"),
  2641 => (x"49",x"72",x"87",x"ce"),
  2642 => (x"c2",x"91",x"cc",x"c1"),
  2643 => (x"c1",x"81",x"f8",x"fb"),
  2644 => (x"79",x"c0",x"81",x"c8"),
  2645 => (x"5e",x"0e",x"4f",x"26"),
  2646 => (x"0e",x"5d",x"5c",x"5b"),
  2647 => (x"4a",x"71",x"86",x"fc"),
  2648 => (x"c0",x"4b",x"d4",x"ff"),
  2649 => (x"4d",x"66",x"d4",x"4c"),
  2650 => (x"01",x"ad",x"b7",x"c3"),
  2651 => (x"72",x"87",x"c2",x"c2"),
  2652 => (x"ec",x"c0",x"02",x"9a"),
  2653 => (x"49",x"75",x"1e",x"87"),
  2654 => (x"c2",x"91",x"cc",x"c1"),
  2655 => (x"71",x"48",x"f8",x"fb"),
  2656 => (x"58",x"a6",x"c8",x"80"),
  2657 => (x"fe",x"49",x"66",x"c4"),
  2658 => (x"c4",x"87",x"fd",x"c2"),
  2659 => (x"02",x"98",x"70",x"86"),
  2660 => (x"49",x"6e",x"87",x"d4"),
  2661 => (x"c1",x"81",x"c8",x"c1"),
  2662 => (x"c8",x"49",x"6e",x"79"),
  2663 => (x"c5",x"4c",x"69",x"81"),
  2664 => (x"fe",x"49",x"75",x"87"),
  2665 => (x"d0",x"ff",x"87",x"d7"),
  2666 => (x"78",x"e1",x"c8",x"48"),
  2667 => (x"48",x"74",x"7b",x"dd"),
  2668 => (x"70",x"98",x"ff",x"c3"),
  2669 => (x"c8",x"49",x"74",x"7b"),
  2670 => (x"48",x"71",x"29",x"b7"),
  2671 => (x"70",x"98",x"ff",x"c3"),
  2672 => (x"d0",x"49",x"74",x"7b"),
  2673 => (x"48",x"71",x"29",x"b7"),
  2674 => (x"70",x"98",x"ff",x"c3"),
  2675 => (x"d8",x"48",x"74",x"7b"),
  2676 => (x"7b",x"70",x"28",x"b7"),
  2677 => (x"7b",x"7b",x"7b",x"c0"),
  2678 => (x"7b",x"7b",x"7b",x"7b"),
  2679 => (x"7b",x"7b",x"7b",x"7b"),
  2680 => (x"48",x"d0",x"ff",x"7b"),
  2681 => (x"75",x"78",x"e0",x"c0"),
  2682 => (x"ff",x"49",x"dc",x"1e"),
  2683 => (x"c4",x"87",x"e6",x"d6"),
  2684 => (x"26",x"8e",x"fc",x"86"),
  2685 => (x"26",x"4c",x"26",x"4d"),
  2686 => (x"14",x"4f",x"26",x"4b"),
  2687 => (x"14",x"00",x"00",x"1d"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

