library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4fec287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49f4fec2",
    18 => x"48cce6c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"c9e6c287",
    25 => x"c5e6c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"edc187f7",
    29 => x"e6c287e6",
    30 => x"e6c24dc9",
    31 => x"ad744cc9",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"5c5b5e0e",
    36 => x"86f00e5d",
    37 => x"a6c44cc0",
    38 => x"c078c048",
    39 => x"c04ba6e4",
    40 => x"484966e0",
    41 => x"e4c080c1",
    42 => x"7e1158a6",
    43 => x"f1c3026e",
    44 => x"0266c487",
    45 => x"c487c6c3",
    46 => x"78c048a6",
    47 => x"f0c04a6e",
    48 => x"dac2028a",
    49 => x"8af3c087",
    50 => x"87dbc202",
    51 => x"dc028ac1",
    52 => x"028ac887",
    53 => x"c487c8c2",
    54 => x"87d1028a",
    55 => x"c1028ac3",
    56 => x"8ac287eb",
    57 => x"c387c602",
    58 => x"c9c2058a",
    59 => x"7383c487",
    60 => x"6989c449",
    61 => x"c1026e7e",
    62 => x"a6c887c8",
    63 => x"c478c048",
    64 => x"cc78c080",
    65 => x"4a6e4d66",
    66 => x"cf2ab7dc",
    67 => x"c4486e9a",
    68 => x"727e7030",
    69 => x"87c5029a",
    70 => x"c148a6c8",
    71 => x"06aac978",
    72 => x"f7c087c5",
    73 => x"c087c382",
    74 => x"66c882f0",
    75 => x"7287c702",
    76 => x"87fac149",
    77 => x"85c184c1",
    78 => x"04adb7c8",
    79 => x"c187c7ff",
    80 => x"f0c087ce",
    81 => x"87e6c149",
    82 => x"c3c184c1",
    83 => x"7383c487",
    84 => x"6a8ac44a",
    85 => x"87f1c149",
    86 => x"4ca44970",
    87 => x"c487f1c0",
    88 => x"78c148a6",
    89 => x"c487e9c0",
    90 => x"c44a7383",
    91 => x"c0496a8a",
    92 => x"84c187fc",
    93 => x"496e87da",
    94 => x"d387f3c0",
    95 => x"c0486e87",
    96 => x"c705a8e5",
    97 => x"48a6c487",
    98 => x"87c478c1",
    99 => x"87de496e",
   100 => x"4966e0c0",
   101 => x"c080c148",
   102 => x"1158a6e4",
   103 => x"fc056e7e",
   104 => x"487487cf",
   105 => x"4d268ef0",
   106 => x"4b264c26",
   107 => x"fc1e4f26",
   108 => x"ff4a7186",
   109 => x"486949c0",
   110 => x"7098c0c4",
   111 => x"0298487e",
   112 => x"797287f4",
   113 => x"268efc48",
   114 => x"5b5e0e4f",
   115 => x"4b710e5c",
   116 => x"4a134cc0",
   117 => x"87cd029a",
   118 => x"d1ff4972",
   119 => x"1384c187",
   120 => x"f3059a4a",
   121 => x"26487487",
   122 => x"264b264c",
   123 => x"1e721e4f",
   124 => x"48121e73",
   125 => x"87ca0211",
   126 => x"98dfc34b",
   127 => x"0288739b",
   128 => x"4b2687f0",
   129 => x"4f264a26",
   130 => x"721e731e",
   131 => x"048bc11e",
   132 => x"481287ca",
   133 => x"87c40211",
   134 => x"87f10288",
   135 => x"4b264a26",
   136 => x"731e4f26",
   137 => x"a9738148",
   138 => x"1287c502",
   139 => x"87f60553",
   140 => x"731e4f26",
   141 => x"c84a711e",
   142 => x"c1494b66",
   143 => x"0299718b",
   144 => x"481287cf",
   145 => x"7808d4ff",
   146 => x"8bc14973",
   147 => x"f1059971",
   148 => x"264b2687",
   149 => x"5b5e0e4f",
   150 => x"4a710e5c",
   151 => x"cc4cd4ff",
   152 => x"c1494b66",
   153 => x"0299718b",
   154 => x"ffc387ce",
   155 => x"73526c7c",
   156 => x"718bc149",
   157 => x"87f20599",
   158 => x"4b264c26",
   159 => x"731e4f26",
   160 => x"4bd4ff1e",
   161 => x"6b7bffc3",
   162 => x"7bffc34a",
   163 => x"32c8496b",
   164 => x"ffc3b172",
   165 => x"c84a6b7b",
   166 => x"c3b27131",
   167 => x"496b7bff",
   168 => x"b17232c8",
   169 => x"4b264871",
   170 => x"5e0e4f26",
   171 => x"0e5d5c5b",
   172 => x"d4ff4d71",
   173 => x"c348754c",
   174 => x"7c7098ff",
   175 => x"bfcce6c2",
   176 => x"d087c805",
   177 => x"30c94866",
   178 => x"d058a6d4",
   179 => x"29d84966",
   180 => x"ffc34871",
   181 => x"d07c7098",
   182 => x"29d04966",
   183 => x"ffc34871",
   184 => x"d07c7098",
   185 => x"29c84966",
   186 => x"ffc34871",
   187 => x"d07c7098",
   188 => x"ffc34866",
   189 => x"757c7098",
   190 => x"7129d049",
   191 => x"98ffc348",
   192 => x"4b6c7c70",
   193 => x"4afff0c9",
   194 => x"05abffc3",
   195 => x"714987cf",
   196 => x"c14b6c7c",
   197 => x"87c5028a",
   198 => x"f202ab71",
   199 => x"26487387",
   200 => x"264c264d",
   201 => x"1e4f264b",
   202 => x"d4ff49c0",
   203 => x"78ffc348",
   204 => x"c8c381c1",
   205 => x"f104a9b7",
   206 => x"0e4f2687",
   207 => x"5d5c5b5e",
   208 => x"f0ffc00e",
   209 => x"c14df7c1",
   210 => x"c0c0c0c0",
   211 => x"d6ff4bc0",
   212 => x"dff8c487",
   213 => x"751ec04c",
   214 => x"87cefd49",
   215 => x"a8c186c4",
   216 => x"87e5c005",
   217 => x"c348d4ff",
   218 => x"1e7378ff",
   219 => x"c1f0e1c0",
   220 => x"f5fc49e9",
   221 => x"7086c487",
   222 => x"87ca0598",
   223 => x"c348d4ff",
   224 => x"48c178ff",
   225 => x"defe87cb",
   226 => x"058cc187",
   227 => x"c087c6ff",
   228 => x"264d2648",
   229 => x"264b264c",
   230 => x"5b5e0e4f",
   231 => x"ffc00e5c",
   232 => x"4cc1c1f0",
   233 => x"c348d4ff",
   234 => x"dccf78ff",
   235 => x"87d9f849",
   236 => x"1ec04bd3",
   237 => x"f1fb4974",
   238 => x"7086c487",
   239 => x"87ca0598",
   240 => x"c348d4ff",
   241 => x"48c178ff",
   242 => x"dafd87cb",
   243 => x"058bc187",
   244 => x"c087dfff",
   245 => x"264c2648",
   246 => x"004f264b",
   247 => x"00444d43",
   248 => x"43484453",
   249 => x"69616620",
   250 => x"000a216c",
   251 => x"52524549",
   252 => x"00000000",
   253 => x"00495053",
   254 => x"74697257",
   255 => x"61662065",
   256 => x"64656c69",
   257 => x"5e0e000a",
   258 => x"0e5d5c5b",
   259 => x"ff4dffc3",
   260 => x"d2fc4bd4",
   261 => x"1eeac687",
   262 => x"c1f0e1c0",
   263 => x"c9fa49c8",
   264 => x"c186c487",
   265 => x"87c802a8",
   266 => x"c087eefd",
   267 => x"87e8c148",
   268 => x"7087cbf9",
   269 => x"ffffcf49",
   270 => x"a9eac699",
   271 => x"fd87c802",
   272 => x"48c087d7",
   273 => x"7587d1c1",
   274 => x"4cf1c07b",
   275 => x"7087ecfb",
   276 => x"ecc00298",
   277 => x"c01ec087",
   278 => x"fac1f0ff",
   279 => x"87caf949",
   280 => x"987086c4",
   281 => x"7587da05",
   282 => x"75496b7b",
   283 => x"757b757b",
   284 => x"c17b757b",
   285 => x"c40299c0",
   286 => x"db48c187",
   287 => x"d748c087",
   288 => x"05acc287",
   289 => x"e0cf87ca",
   290 => x"87fdf449",
   291 => x"87c848c0",
   292 => x"fe058cc1",
   293 => x"48c087f6",
   294 => x"4c264d26",
   295 => x"4f264b26",
   296 => x"5c5b5e0e",
   297 => x"d0ff0e5d",
   298 => x"d0e5c04d",
   299 => x"c24cc0c1",
   300 => x"c148cce6",
   301 => x"49f4cf78",
   302 => x"c787cef4",
   303 => x"f97dc24b",
   304 => x"7dc387e5",
   305 => x"49741ec0",
   306 => x"c487dff7",
   307 => x"05a8c186",
   308 => x"c24b87c1",
   309 => x"87cb05ab",
   310 => x"f349eccf",
   311 => x"48c087eb",
   312 => x"c187f6c0",
   313 => x"d4ff058b",
   314 => x"87dafc87",
   315 => x"58d0e6c2",
   316 => x"cd059870",
   317 => x"c01ec187",
   318 => x"d0c1f0ff",
   319 => x"87eaf649",
   320 => x"d4ff86c4",
   321 => x"78ffc348",
   322 => x"c287eec4",
   323 => x"c258d4e6",
   324 => x"48d4ff7d",
   325 => x"c178ffc3",
   326 => x"264d2648",
   327 => x"264b264c",
   328 => x"5b5e0e4f",
   329 => x"710e5d5c",
   330 => x"4cffc34d",
   331 => x"744bd4ff",
   332 => x"48d0ff7b",
   333 => x"7478c3c4",
   334 => x"c01e757b",
   335 => x"d8c1f0ff",
   336 => x"87e6f549",
   337 => x"987086c4",
   338 => x"cf87cb02",
   339 => x"f8f149f8",
   340 => x"c048c187",
   341 => x"7b7487ee",
   342 => x"c87bfec3",
   343 => x"66d41ec0",
   344 => x"87cef349",
   345 => x"7b7486c4",
   346 => x"7b747b74",
   347 => x"4ae0dad8",
   348 => x"056b7b74",
   349 => x"8ac187c5",
   350 => x"7487f505",
   351 => x"48d0ff7b",
   352 => x"48c078c2",
   353 => x"4c264d26",
   354 => x"4f264b26",
   355 => x"5c5b5e0e",
   356 => x"86fc0e5d",
   357 => x"d4ff4b71",
   358 => x"c57ec04c",
   359 => x"4adfcdee",
   360 => x"6c7cffc3",
   361 => x"a8fec348",
   362 => x"87f8c005",
   363 => x"9b734d74",
   364 => x"d487cc02",
   365 => x"49731e66",
   366 => x"c487daf2",
   367 => x"ff87d486",
   368 => x"d1c448d0",
   369 => x"4a66d478",
   370 => x"c17dffc3",
   371 => x"87f8058a",
   372 => x"c35aa6d8",
   373 => x"737c7cff",
   374 => x"87c5059b",
   375 => x"d048d0ff",
   376 => x"7e4ac178",
   377 => x"fe058ac1",
   378 => x"486e87f6",
   379 => x"4d268efc",
   380 => x"4b264c26",
   381 => x"731e4f26",
   382 => x"c04a711e",
   383 => x"48d4ff4b",
   384 => x"ff78ffc3",
   385 => x"c3c448d0",
   386 => x"48d4ff78",
   387 => x"7278ffc3",
   388 => x"f0ffc01e",
   389 => x"f249d1c1",
   390 => x"86c487d0",
   391 => x"d2059870",
   392 => x"1ec0c887",
   393 => x"fd4966cc",
   394 => x"86c487e2",
   395 => x"d0ff4b70",
   396 => x"7378c248",
   397 => x"264b2648",
   398 => x"5b5e0e4f",
   399 => x"c00e5d5c",
   400 => x"f0ffc01e",
   401 => x"f149c9c1",
   402 => x"1ed287e0",
   403 => x"49dce6c2",
   404 => x"c887f9fc",
   405 => x"c14cc086",
   406 => x"acb7d284",
   407 => x"c287f804",
   408 => x"bf97dce6",
   409 => x"99c0c349",
   410 => x"05a9c0c1",
   411 => x"c287e7c0",
   412 => x"bf97e3e6",
   413 => x"c231d049",
   414 => x"bf97e4e6",
   415 => x"7232c84a",
   416 => x"e5e6c2b1",
   417 => x"b14abf97",
   418 => x"ffcf4c71",
   419 => x"c19cffff",
   420 => x"c134ca84",
   421 => x"e6c287e7",
   422 => x"49bf97e5",
   423 => x"99c631c1",
   424 => x"97e6e6c2",
   425 => x"b7c74abf",
   426 => x"c2b1722a",
   427 => x"bf97e1e6",
   428 => x"9dcf4d4a",
   429 => x"97e2e6c2",
   430 => x"9ac34abf",
   431 => x"e6c232ca",
   432 => x"4bbf97e3",
   433 => x"b27333c2",
   434 => x"97e4e6c2",
   435 => x"c0c34bbf",
   436 => x"2bb7c69b",
   437 => x"81c2b273",
   438 => x"307148c1",
   439 => x"48c14970",
   440 => x"4d703075",
   441 => x"84c14c72",
   442 => x"c0c89471",
   443 => x"cc06adb7",
   444 => x"b734c187",
   445 => x"b7c0c82d",
   446 => x"f4ff01ad",
   447 => x"26487487",
   448 => x"264c264d",
   449 => x"0e4f264b",
   450 => x"5d5c5b5e",
   451 => x"c286fc0e",
   452 => x"c048c4ef",
   453 => x"fce6c278",
   454 => x"fb49c01e",
   455 => x"86c487d8",
   456 => x"c5059870",
   457 => x"c948c087",
   458 => x"4dc087d5",
   459 => x"48c0f4c2",
   460 => x"e7c278c1",
   461 => x"e6c04af2",
   462 => x"4bc849d8",
   463 => x"7087c9eb",
   464 => x"87c60598",
   465 => x"48c0f4c2",
   466 => x"e8c278c0",
   467 => x"e6c04ace",
   468 => x"4bc849e4",
   469 => x"7087f1ea",
   470 => x"87c60598",
   471 => x"48c0f4c2",
   472 => x"f4c278c0",
   473 => x"c002bfc0",
   474 => x"eec287fe",
   475 => x"c24dbfc2",
   476 => x"bf9ffaee",
   477 => x"c5486e7e",
   478 => x"05a8ead6",
   479 => x"eec287c7",
   480 => x"ce4dbfc2",
   481 => x"ca486e87",
   482 => x"02a8d5e9",
   483 => x"48c087c5",
   484 => x"c287ecc7",
   485 => x"751efce6",
   486 => x"87daf949",
   487 => x"987086c4",
   488 => x"c087c505",
   489 => x"87d7c748",
   490 => x"4acee8c2",
   491 => x"49f0e6c0",
   492 => x"d3e94bc8",
   493 => x"05987087",
   494 => x"c287c8c0",
   495 => x"c148c4ef",
   496 => x"c287d878",
   497 => x"c04af2e7",
   498 => x"c849fce6",
   499 => x"87f8e84b",
   500 => x"c0029870",
   501 => x"48c087c5",
   502 => x"c287e4c6",
   503 => x"bf97faee",
   504 => x"a9d5c149",
   505 => x"87cdc005",
   506 => x"97fbeec2",
   507 => x"eac249bf",
   508 => x"c5c002a9",
   509 => x"c648c087",
   510 => x"e6c287c5",
   511 => x"7ebf97fc",
   512 => x"e9c3486e",
   513 => x"cec002a8",
   514 => x"c3486e87",
   515 => x"c002a8eb",
   516 => x"48c087c5",
   517 => x"c287e8c5",
   518 => x"bf97c7e7",
   519 => x"c0059949",
   520 => x"e7c287cc",
   521 => x"49bf97c8",
   522 => x"c002a9c2",
   523 => x"48c087c5",
   524 => x"c287ccc5",
   525 => x"bf97c9e7",
   526 => x"c0efc248",
   527 => x"484c7058",
   528 => x"efc288c1",
   529 => x"e7c258c4",
   530 => x"49bf97ca",
   531 => x"e7c28175",
   532 => x"4abf97cb",
   533 => x"a17232c8",
   534 => x"dcf3c27e",
   535 => x"c2786e48",
   536 => x"bf97cce7",
   537 => x"f4f3c248",
   538 => x"c4efc258",
   539 => x"d3c202bf",
   540 => x"cee8c287",
   541 => x"cce6c04a",
   542 => x"e64bc849",
   543 => x"987087ca",
   544 => x"87c5c002",
   545 => x"f6c348c0",
   546 => x"fceec287",
   547 => x"f3c24cbf",
   548 => x"e7c25cf0",
   549 => x"49bf97e1",
   550 => x"e7c231c8",
   551 => x"4abf97e0",
   552 => x"e7c249a1",
   553 => x"4abf97e2",
   554 => x"a17232d0",
   555 => x"e3e7c249",
   556 => x"d84abf97",
   557 => x"49a17232",
   558 => x"59f8f3c2",
   559 => x"bff0f3c2",
   560 => x"dcf3c291",
   561 => x"f3c281bf",
   562 => x"e7c259e4",
   563 => x"4abf97e9",
   564 => x"e7c232c8",
   565 => x"4bbf97e8",
   566 => x"e7c24aa2",
   567 => x"4bbf97ea",
   568 => x"a27333d0",
   569 => x"ebe7c24a",
   570 => x"cf4bbf97",
   571 => x"7333d89b",
   572 => x"f3c24aa2",
   573 => x"8ac25ae8",
   574 => x"f3c29274",
   575 => x"a17248e8",
   576 => x"87c7c178",
   577 => x"97cee7c2",
   578 => x"31c849bf",
   579 => x"97cde7c2",
   580 => x"49a14abf",
   581 => x"ffc731c5",
   582 => x"c229c981",
   583 => x"c259f0f3",
   584 => x"bf97d3e7",
   585 => x"c232c84a",
   586 => x"bf97d2e7",
   587 => x"c24aa24b",
   588 => x"c25af8f3",
   589 => x"92bff0f3",
   590 => x"f3c2826e",
   591 => x"f3c25aec",
   592 => x"78c048e4",
   593 => x"48e0f3c2",
   594 => x"c278a172",
   595 => x"c248f8f3",
   596 => x"78bfe4f3",
   597 => x"48fcf3c2",
   598 => x"bfe8f3c2",
   599 => x"c4efc278",
   600 => x"c9c002bf",
   601 => x"c4487487",
   602 => x"c07e7030",
   603 => x"f3c287c9",
   604 => x"c448bfec",
   605 => x"c27e7030",
   606 => x"6e48c8ef",
   607 => x"fc48c178",
   608 => x"264d268e",
   609 => x"264b264c",
   610 => x"0000004f",
   611 => x"33544146",
   612 => x"20202032",
   613 => x"00000000",
   614 => x"31544146",
   615 => x"20202036",
   616 => x"00000000",
   617 => x"33544146",
   618 => x"20202032",
   619 => x"00000000",
   620 => x"33544146",
   621 => x"20202032",
   622 => x"00000000",
   623 => x"31544146",
   624 => x"20202036",
   625 => x"5b5e0e00",
   626 => x"710e5d5c",
   627 => x"c4efc24a",
   628 => x"87cb02bf",
   629 => x"2bc74b72",
   630 => x"ffc14d72",
   631 => x"7287c99d",
   632 => x"722bc84b",
   633 => x"9dffc34d",
   634 => x"bfdcf3c2",
   635 => x"d0fec083",
   636 => x"d902abbf",
   637 => x"d4fec087",
   638 => x"fce6c25b",
   639 => x"ef49731e",
   640 => x"86c487f4",
   641 => x"c5059870",
   642 => x"c048c087",
   643 => x"efc287e6",
   644 => x"d202bfc4",
   645 => x"c4497587",
   646 => x"fce6c291",
   647 => x"cf4c6981",
   648 => x"ffffffff",
   649 => x"7587cb9c",
   650 => x"c291c249",
   651 => x"9f81fce6",
   652 => x"48744c69",
   653 => x"4c264d26",
   654 => x"4f264b26",
   655 => x"5c5b5e0e",
   656 => x"86f40e5d",
   657 => x"c459a6c8",
   658 => x"80c84866",
   659 => x"486e7e70",
   660 => x"c11e78c0",
   661 => x"87fdcc49",
   662 => x"4c7086c4",
   663 => x"fcc0029c",
   664 => x"ccefc287",
   665 => x"4966dc4a",
   666 => x"87c1deff",
   667 => x"c0029870",
   668 => x"4a7487eb",
   669 => x"cb4966dc",
   670 => x"cbdeff4b",
   671 => x"02987087",
   672 => x"1ec087db",
   673 => x"c4029c74",
   674 => x"c24dc087",
   675 => x"754dc187",
   676 => x"87c1cc49",
   677 => x"4c7086c4",
   678 => x"c4ff059c",
   679 => x"029c7487",
   680 => x"dc87f4c1",
   681 => x"486e49a4",
   682 => x"a4da7869",
   683 => x"4d66c449",
   684 => x"699f85c4",
   685 => x"c4efc27d",
   686 => x"87d202bf",
   687 => x"9f49a4d4",
   688 => x"ffc04969",
   689 => x"487199ff",
   690 => x"7e7030d0",
   691 => x"7ec087c2",
   692 => x"6d48496e",
   693 => x"c47d7080",
   694 => x"78c04866",
   695 => x"cc4966c4",
   696 => x"c4796d81",
   697 => x"81d04966",
   698 => x"a6c879c0",
   699 => x"c878c048",
   700 => x"66c44c66",
   701 => x"7482d44a",
   702 => x"7291c849",
   703 => x"41c049a1",
   704 => x"84c1796d",
   705 => x"04acb7c6",
   706 => x"c487e7ff",
   707 => x"c4c14966",
   708 => x"c179c081",
   709 => x"c087c248",
   710 => x"268ef448",
   711 => x"264c264d",
   712 => x"0e4f264b",
   713 => x"5d5c5b5e",
   714 => x"d04c710e",
   715 => x"496c4d66",
   716 => x"c2b97585",
   717 => x"4abfc0ef",
   718 => x"9972baff",
   719 => x"c0029971",
   720 => x"a4c487e4",
   721 => x"f9496b4b",
   722 => x"7b7087fb",
   723 => x"bffceec2",
   724 => x"71816c49",
   725 => x"c2b9757c",
   726 => x"4abfc0ef",
   727 => x"9972baff",
   728 => x"ff059971",
   729 => x"7c7587dc",
   730 => x"4c264d26",
   731 => x"4f264b26",
   732 => x"711e731e",
   733 => x"e0f3c24b",
   734 => x"a3c449bf",
   735 => x"c24a6a4a",
   736 => x"fceec28a",
   737 => x"a17292bf",
   738 => x"c0efc249",
   739 => x"9a6b4abf",
   740 => x"c049a172",
   741 => x"c859d4fe",
   742 => x"e9711e66",
   743 => x"86c487d8",
   744 => x"c4059870",
   745 => x"c248c087",
   746 => x"2648c187",
   747 => x"1e4f264b",
   748 => x"4b711e73",
   749 => x"bfe0f3c2",
   750 => x"4aa3c449",
   751 => x"8ac24a6a",
   752 => x"bffceec2",
   753 => x"49a17292",
   754 => x"bfc0efc2",
   755 => x"729a6b4a",
   756 => x"fec049a1",
   757 => x"66c859d4",
   758 => x"c4e5711e",
   759 => x"7086c487",
   760 => x"87c40598",
   761 => x"87c248c0",
   762 => x"4b2648c1",
   763 => x"5e0e4f26",
   764 => x"0e5d5c5b",
   765 => x"4b7186e4",
   766 => x"4866ecc0",
   767 => x"a6cc28c9",
   768 => x"c0efc258",
   769 => x"b9ff49bf",
   770 => x"66c84871",
   771 => x"58a6d498",
   772 => x"986b4871",
   773 => x"c458a6d0",
   774 => x"a6c47ea3",
   775 => x"78bf6e48",
   776 => x"cc4866d0",
   777 => x"c605a866",
   778 => x"7b66c887",
   779 => x"d487c6c3",
   780 => x"ffc148a6",
   781 => x"ffffffff",
   782 => x"ff80c478",
   783 => x"d44ac078",
   784 => x"49724da3",
   785 => x"a17591c8",
   786 => x"4c66d049",
   787 => x"b7c08c69",
   788 => x"87cd04ac",
   789 => x"acb766d4",
   790 => x"dc87c603",
   791 => x"a6d85aa6",
   792 => x"c682c15c",
   793 => x"ff04aab7",
   794 => x"66d887d5",
   795 => x"a8b7c048",
   796 => x"d887d004",
   797 => x"91c84966",
   798 => x"2149a175",
   799 => x"69486e7b",
   800 => x"c087c978",
   801 => x"49a3cc7b",
   802 => x"7869486e",
   803 => x"6b4866c8",
   804 => x"58a6cc88",
   805 => x"bffceec2",
   806 => x"7090c848",
   807 => x"4866c87e",
   808 => x"c901a86e",
   809 => x"4866c887",
   810 => x"c003a86e",
   811 => x"c4c187fd",
   812 => x"bf6e7ea3",
   813 => x"7591c849",
   814 => x"66cc49a1",
   815 => x"49bf6e79",
   816 => x"a17591c8",
   817 => x"6681c449",
   818 => x"48a6d079",
   819 => x"d078bf6e",
   820 => x"a8c54866",
   821 => x"c487c705",
   822 => x"78c048a6",
   823 => x"66d087c8",
   824 => x"c880c148",
   825 => x"486e58a6",
   826 => x"c87866c4",
   827 => x"49731e66",
   828 => x"c487f0f8",
   829 => x"fce6c286",
   830 => x"f949731e",
   831 => x"a3d087f2",
   832 => x"66f0c049",
   833 => x"268ee079",
   834 => x"264c264d",
   835 => x"0e4f264b",
   836 => x"0e5c5b5e",
   837 => x"4bc04a71",
   838 => x"c0029a72",
   839 => x"a2da87e0",
   840 => x"4b699f49",
   841 => x"bfc4efc2",
   842 => x"d487cf02",
   843 => x"699f49a2",
   844 => x"ffc04c49",
   845 => x"34d09cff",
   846 => x"4cc087c2",
   847 => x"9b73b374",
   848 => x"4a87df02",
   849 => x"eec28ac2",
   850 => x"9249bffc",
   851 => x"bfe0f3c2",
   852 => x"c2807248",
   853 => x"7158c0f4",
   854 => x"c230c448",
   855 => x"c058ccef",
   856 => x"f3c287e9",
   857 => x"c24bbfe4",
   858 => x"c248fcf3",
   859 => x"78bfe8f3",
   860 => x"bfc4efc2",
   861 => x"c287c902",
   862 => x"49bffcee",
   863 => x"87c731c4",
   864 => x"bfecf3c2",
   865 => x"c231c449",
   866 => x"c259ccef",
   867 => x"265bfcf3",
   868 => x"264b264c",
   869 => x"5b5e0e4f",
   870 => x"f00e5d5c",
   871 => x"59a6c886",
   872 => x"ffffffcf",
   873 => x"7ec04cf8",
   874 => x"d80266c4",
   875 => x"f8e6c287",
   876 => x"c278c048",
   877 => x"c248f0e6",
   878 => x"78bffcf3",
   879 => x"48f4e6c2",
   880 => x"bff8f3c2",
   881 => x"d9efc278",
   882 => x"c250c048",
   883 => x"49bfc8ef",
   884 => x"bff8e6c2",
   885 => x"03aa714a",
   886 => x"7287ccc4",
   887 => x"0599cf49",
   888 => x"c087eac0",
   889 => x"c248d0fe",
   890 => x"78bff0e6",
   891 => x"1efce6c2",
   892 => x"bff0e6c2",
   893 => x"f0e6c249",
   894 => x"78a1c148",
   895 => x"f5dfff71",
   896 => x"c086c487",
   897 => x"c248ccfe",
   898 => x"cc78fce6",
   899 => x"ccfec087",
   900 => x"e0c048bf",
   901 => x"d0fec080",
   902 => x"f8e6c258",
   903 => x"80c148bf",
   904 => x"58fce6c2",
   905 => x"000f8c27",
   906 => x"bf97bf00",
   907 => x"c2029d4d",
   908 => x"e5c387e5",
   909 => x"dec202ad",
   910 => x"ccfec087",
   911 => x"a3cb4bbf",
   912 => x"cf4c1149",
   913 => x"d2c105ac",
   914 => x"df497587",
   915 => x"cd89c199",
   916 => x"ccefc291",
   917 => x"4aa3c181",
   918 => x"a3c35112",
   919 => x"c551124a",
   920 => x"51124aa3",
   921 => x"124aa3c7",
   922 => x"4aa3c951",
   923 => x"a3ce5112",
   924 => x"d051124a",
   925 => x"51124aa3",
   926 => x"124aa3d2",
   927 => x"4aa3d451",
   928 => x"a3d65112",
   929 => x"d851124a",
   930 => x"51124aa3",
   931 => x"124aa3dc",
   932 => x"4aa3de51",
   933 => x"7ec15112",
   934 => x"7487fcc0",
   935 => x"0599c849",
   936 => x"7487edc0",
   937 => x"0599d049",
   938 => x"e0c087d3",
   939 => x"ccc00266",
   940 => x"c0497387",
   941 => x"700f66e0",
   942 => x"d3c00298",
   943 => x"c0056e87",
   944 => x"efc287c6",
   945 => x"50c048cc",
   946 => x"bfccfec0",
   947 => x"87e9c248",
   948 => x"48d9efc2",
   949 => x"c27e50c0",
   950 => x"49bfc8ef",
   951 => x"bff8e6c2",
   952 => x"04aa714a",
   953 => x"cf87f4fb",
   954 => x"f8ffffff",
   955 => x"fcf3c24c",
   956 => x"c8c005bf",
   957 => x"c4efc287",
   958 => x"fac102bf",
   959 => x"f4e6c287",
   960 => x"c0eb49bf",
   961 => x"f8e6c287",
   962 => x"48a6c458",
   963 => x"bff4e6c2",
   964 => x"c4efc278",
   965 => x"dbc002bf",
   966 => x"4966c487",
   967 => x"a9749974",
   968 => x"87c8c002",
   969 => x"c048a6c8",
   970 => x"87e7c078",
   971 => x"c148a6c8",
   972 => x"87dfc078",
   973 => x"cf4966c4",
   974 => x"a999f8ff",
   975 => x"87c8c002",
   976 => x"c048a6cc",
   977 => x"87c5c078",
   978 => x"c148a6cc",
   979 => x"48a6c878",
   980 => x"c87866cc",
   981 => x"dec00566",
   982 => x"4966c487",
   983 => x"eec289c2",
   984 => x"c291bffc",
   985 => x"48bfe0f3",
   986 => x"e6c28071",
   987 => x"e6c258f4",
   988 => x"78c048f8",
   989 => x"c087d4f9",
   990 => x"ffffcf48",
   991 => x"f04cf8ff",
   992 => x"264d268e",
   993 => x"264b264c",
   994 => x"0000004f",
   995 => x"00000000",
   996 => x"ffffffff",
   997 => x"48d4ff1e",
   998 => x"2678ffc3",
   999 => x"d4ff1e4f",
  1000 => x"78ffc348",
  1001 => x"c048d0ff",
  1002 => x"d4ff78e1",
  1003 => x"2678d448",
  1004 => x"d0ff1e4f",
  1005 => x"78e0c048",
  1006 => x"ff1e4f26",
  1007 => x"497087d6",
  1008 => x"87c60299",
  1009 => x"05a9fbc0",
  1010 => x"487187f1",
  1011 => x"5e0e4f26",
  1012 => x"710e5c5b",
  1013 => x"fe4cc04b",
  1014 => x"497087fa",
  1015 => x"f9c00299",
  1016 => x"a9ecc087",
  1017 => x"87f2c002",
  1018 => x"02a9fbc0",
  1019 => x"cc87ebc0",
  1020 => x"03acb766",
  1021 => x"66d087c7",
  1022 => x"7187c202",
  1023 => x"02997153",
  1024 => x"84c187c2",
  1025 => x"7087cdfe",
  1026 => x"cd029949",
  1027 => x"a9ecc087",
  1028 => x"c087c702",
  1029 => x"ff05a9fb",
  1030 => x"66d087d5",
  1031 => x"c087c302",
  1032 => x"fbc07b97",
  1033 => x"87c705a9",
  1034 => x"0ac04a74",
  1035 => x"7487c28a",
  1036 => x"2648724a",
  1037 => x"264b264c",
  1038 => x"d7fd1e4f",
  1039 => x"c0497087",
  1040 => x"c904a9f0",
  1041 => x"a9f9c087",
  1042 => x"c087c301",
  1043 => x"c1c189f0",
  1044 => x"87c904a9",
  1045 => x"01a9dac1",
  1046 => x"f7c087c3",
  1047 => x"26487189",
  1048 => x"5b5e0e4f",
  1049 => x"f80e5d5c",
  1050 => x"c04c7186",
  1051 => x"87edfc7e",
  1052 => x"c4c14bc0",
  1053 => x"49bf97c0",
  1054 => x"cf04a9c0",
  1055 => x"87fafc87",
  1056 => x"c4c183c1",
  1057 => x"49bf97c0",
  1058 => x"87f106ab",
  1059 => x"97c0c4c1",
  1060 => x"87cf02bf",
  1061 => x"7087fdfb",
  1062 => x"c6029949",
  1063 => x"a9ecc087",
  1064 => x"c087f105",
  1065 => x"87ecfb4b",
  1066 => x"e7fb4d70",
  1067 => x"58a6c887",
  1068 => x"7087e1fb",
  1069 => x"c883c14a",
  1070 => x"699749a4",
  1071 => x"da05ad49",
  1072 => x"49a4c987",
  1073 => x"c4496997",
  1074 => x"ce05a966",
  1075 => x"49a4ca87",
  1076 => x"aa496997",
  1077 => x"c187c405",
  1078 => x"c087d07e",
  1079 => x"c602adec",
  1080 => x"adfbc087",
  1081 => x"c087c405",
  1082 => x"6e7ec14b",
  1083 => x"87f5fe02",
  1084 => x"7387fefa",
  1085 => x"268ef848",
  1086 => x"264c264d",
  1087 => x"004f264b",
  1088 => x"1e731e00",
  1089 => x"c84bd4ff",
  1090 => x"d0ff4a66",
  1091 => x"78c5c848",
  1092 => x"c148d4ff",
  1093 => x"7b1178d4",
  1094 => x"f9058ac1",
  1095 => x"48d0ff87",
  1096 => x"4b2678c4",
  1097 => x"5e0e4f26",
  1098 => x"0e5d5c5b",
  1099 => x"7e7186f8",
  1100 => x"f4c21e6e",
  1101 => x"c3e449d0",
  1102 => x"7086c487",
  1103 => x"edc40298",
  1104 => x"dcf1c187",
  1105 => x"496e4cbf",
  1106 => x"c887d6fc",
  1107 => x"c9c158a6",
  1108 => x"fcfe1efc",
  1109 => x"86c487f6",
  1110 => x"87c50566",
  1111 => x"c148a6c4",
  1112 => x"48d0ff78",
  1113 => x"d4ff78c5",
  1114 => x"78d5c148",
  1115 => x"c14966c4",
  1116 => x"c131c689",
  1117 => x"bf97d4f1",
  1118 => x"b071484a",
  1119 => x"7808d4ff",
  1120 => x"c448d0ff",
  1121 => x"ccf4c278",
  1122 => x"d049bf97",
  1123 => x"87dd0299",
  1124 => x"d4ff78c5",
  1125 => x"78d6c148",
  1126 => x"d4ff4ac0",
  1127 => x"78ffc348",
  1128 => x"e0c082c1",
  1129 => x"87f204aa",
  1130 => x"c448d0ff",
  1131 => x"48d4ff78",
  1132 => x"ff78ffc3",
  1133 => x"78c548d0",
  1134 => x"c148d4ff",
  1135 => x"78c178d3",
  1136 => x"c448d0ff",
  1137 => x"acb7c078",
  1138 => x"87cbc206",
  1139 => x"bfd8f4c2",
  1140 => x"7e748c4b",
  1141 => x"c1029b73",
  1142 => x"c0c887dd",
  1143 => x"b7c08b4d",
  1144 => x"87c603ab",
  1145 => x"4da3c0c8",
  1146 => x"f4c24bc0",
  1147 => x"49bf97cc",
  1148 => x"cf0299d0",
  1149 => x"c21ec087",
  1150 => x"e549d0f4",
  1151 => x"86c487f2",
  1152 => x"87d84c70",
  1153 => x"1efce6c2",
  1154 => x"49d0f4c2",
  1155 => x"7087e1e5",
  1156 => x"c21e754c",
  1157 => x"fb49fce6",
  1158 => x"86c887e7",
  1159 => x"c5059c74",
  1160 => x"c148c087",
  1161 => x"1ec187ca",
  1162 => x"49d0f4c2",
  1163 => x"c487f4e3",
  1164 => x"059b7386",
  1165 => x"6e87e3fe",
  1166 => x"acb7c04c",
  1167 => x"c287d106",
  1168 => x"c048d0f4",
  1169 => x"c080d078",
  1170 => x"c280f478",
  1171 => x"78bfdcf4",
  1172 => x"01acb7c0",
  1173 => x"ff87f5fd",
  1174 => x"78c548d0",
  1175 => x"c148d4ff",
  1176 => x"78c078d3",
  1177 => x"c448d0ff",
  1178 => x"c048c178",
  1179 => x"48c087c2",
  1180 => x"4d268ef8",
  1181 => x"4b264c26",
  1182 => x"00004f26",
  1183 => x"20746f47",
  1184 => x"69747865",
  1185 => x"0000646e",
  1186 => x"64616f4c",
  1187 => x"2e676e69",
  1188 => x"00002e2e",
  1189 => x"61422080",
  1190 => x"00006b63",
  1191 => x"64616f4c",
  1192 => x"202e2a20",
  1193 => x"00000000",
  1194 => x"0000203a",
  1195 => x"61422080",
  1196 => x"00006b63",
  1197 => x"78452080",
  1198 => x"00007469",
  1199 => x"49204453",
  1200 => x"2e74696e",
  1201 => x"0000002e",
  1202 => x"00004b4f",
  1203 => x"544f4f42",
  1204 => x"20202020",
  1205 => x"004d4f52",
  1206 => x"5c5b5e0e",
  1207 => x"86fc0e5d",
  1208 => x"4bc04d71",
  1209 => x"c004ad4c",
  1210 => x"c1c187e8",
  1211 => x"9c741ee1",
  1212 => x"c087c402",
  1213 => x"c187c24a",
  1214 => x"ea49724a",
  1215 => x"86c487d7",
  1216 => x"83c17e70",
  1217 => x"87c2056e",
  1218 => x"84c14b75",
  1219 => x"ff06ab75",
  1220 => x"486e87d8",
  1221 => x"4d268efc",
  1222 => x"4b264c26",
  1223 => x"5e0e4f26",
  1224 => x"0e5d5c5b",
  1225 => x"4d7186f4",
  1226 => x"c291de49",
  1227 => x"7148f0f5",
  1228 => x"6e7e7080",
  1229 => x"c202bf97",
  1230 => x"f5c287cb",
  1231 => x"7549bfe0",
  1232 => x"d3fe7181",
  1233 => x"58a6c887",
  1234 => x"c10266c4",
  1235 => x"f5c287e1",
  1236 => x"66c44be4",
  1237 => x"fe49cb4a",
  1238 => x"7587c7fb",
  1239 => x"c193cc4b",
  1240 => x"c483e0f1",
  1241 => x"c8cac183",
  1242 => x"c149757b",
  1243 => x"6e87fdc0",
  1244 => x"d8f1c17b",
  1245 => x"cc48bf97",
  1246 => x"987058a6",
  1247 => x"4887db02",
  1248 => x"7088f0c0",
  1249 => x"0298487e",
  1250 => x"c14c87d9",
  1251 => x"87d3028c",
  1252 => x"87cf028c",
  1253 => x"87cb028c",
  1254 => x"f5c287d5",
  1255 => x"c5f649e4",
  1256 => x"6e87cc87",
  1257 => x"e4f5c21e",
  1258 => x"f3d4c149",
  1259 => x"7586c487",
  1260 => x"f7ffc049",
  1261 => x"c149c087",
  1262 => x"c287d2c1",
  1263 => x"c048c8f4",
  1264 => x"e2df4950",
  1265 => x"268ef487",
  1266 => x"264c264d",
  1267 => x"1e4f264b",
  1268 => x"4b711e73",
  1269 => x"e0f5c249",
  1270 => x"fb7181bf",
  1271 => x"4a7087fa",
  1272 => x"87c4029a",
  1273 => x"87e7e449",
  1274 => x"48e0f5c2",
  1275 => x"497378c0",
  1276 => x"2687fac1",
  1277 => x"1e4f264b",
  1278 => x"4b711e73",
  1279 => x"024aa3c4",
  1280 => x"c187d0c1",
  1281 => x"87dc028a",
  1282 => x"f2c0028a",
  1283 => x"c1058a87",
  1284 => x"f5c287d3",
  1285 => x"c102bfe0",
  1286 => x"c14887cb",
  1287 => x"e4f5c288",
  1288 => x"87c1c158",
  1289 => x"bfe0f5c2",
  1290 => x"c289c649",
  1291 => x"c059e4f5",
  1292 => x"c003a9b7",
  1293 => x"f5c287ef",
  1294 => x"78c048e0",
  1295 => x"c287e6c0",
  1296 => x"02bfdcf5",
  1297 => x"f5c287df",
  1298 => x"c148bfe0",
  1299 => x"e4f5c280",
  1300 => x"c287d258",
  1301 => x"02bfdcf5",
  1302 => x"f5c287cb",
  1303 => x"c648bfe0",
  1304 => x"e4f5c280",
  1305 => x"c4497358",
  1306 => x"264b2687",
  1307 => x"5b5e0e4f",
  1308 => x"f00e5d5c",
  1309 => x"59a6d086",
  1310 => x"4dfce6c2",
  1311 => x"f5c24cc0",
  1312 => x"78c148dc",
  1313 => x"c048a6c8",
  1314 => x"c27e7578",
  1315 => x"48bfe0f5",
  1316 => x"c106a8c0",
  1317 => x"a6c887c0",
  1318 => x"c27e755c",
  1319 => x"9848fce6",
  1320 => x"87f2c002",
  1321 => x"c14d66c4",
  1322 => x"cc1ee1c1",
  1323 => x"87c40266",
  1324 => x"87c24cc0",
  1325 => x"49744cc1",
  1326 => x"c487dae3",
  1327 => x"c17e7086",
  1328 => x"4866c885",
  1329 => x"a6cc80c1",
  1330 => x"e0f5c258",
  1331 => x"c503adbf",
  1332 => x"ff056e87",
  1333 => x"4d6e87d1",
  1334 => x"9d754cc0",
  1335 => x"87dcc302",
  1336 => x"1ee1c1c1",
  1337 => x"c70266cc",
  1338 => x"48a6c887",
  1339 => x"87c578c0",
  1340 => x"c148a6c8",
  1341 => x"4966c878",
  1342 => x"c487dae2",
  1343 => x"487e7086",
  1344 => x"e4c20298",
  1345 => x"81cb4987",
  1346 => x"d0496997",
  1347 => x"d4c10299",
  1348 => x"cc497487",
  1349 => x"e0f1c191",
  1350 => x"cfcfc181",
  1351 => x"c381c879",
  1352 => x"497451ff",
  1353 => x"f5c291de",
  1354 => x"85714df0",
  1355 => x"7d97c1c2",
  1356 => x"c049a5c1",
  1357 => x"efc251e0",
  1358 => x"02bf97cc",
  1359 => x"84c187d2",
  1360 => x"c24ba5c2",
  1361 => x"db4accef",
  1362 => x"d5f3fe49",
  1363 => x"87d9c187",
  1364 => x"c049a5cd",
  1365 => x"c284c151",
  1366 => x"4a6e4ba5",
  1367 => x"f3fe49cb",
  1368 => x"c4c187c0",
  1369 => x"cc497487",
  1370 => x"e0f1c191",
  1371 => x"deccc181",
  1372 => x"ccefc279",
  1373 => x"d802bf97",
  1374 => x"de497487",
  1375 => x"c284c191",
  1376 => x"714bf0f5",
  1377 => x"ccefc283",
  1378 => x"fe49dd4a",
  1379 => x"d887d3f2",
  1380 => x"de4b7487",
  1381 => x"f0f5c293",
  1382 => x"49a3cb83",
  1383 => x"84c151c0",
  1384 => x"cb4a6e73",
  1385 => x"f9f1fe49",
  1386 => x"4866c887",
  1387 => x"a6cc80c1",
  1388 => x"03acc758",
  1389 => x"6e87c5c0",
  1390 => x"87e4fc05",
  1391 => x"c003acc7",
  1392 => x"f5c287e4",
  1393 => x"78c048dc",
  1394 => x"91cc4974",
  1395 => x"81e0f1c1",
  1396 => x"79deccc1",
  1397 => x"91de4974",
  1398 => x"81f0f5c2",
  1399 => x"84c151c0",
  1400 => x"ff04acc7",
  1401 => x"f2c187dc",
  1402 => x"50c048fc",
  1403 => x"d9c180f7",
  1404 => x"cac140c5",
  1405 => x"80c878d4",
  1406 => x"78f7cfc1",
  1407 => x"c04966cc",
  1408 => x"f087e9f6",
  1409 => x"264d268e",
  1410 => x"264b264c",
  1411 => x"1e731e4f",
  1412 => x"cc494b71",
  1413 => x"e0f1c191",
  1414 => x"4aa1c881",
  1415 => x"48d4f1c1",
  1416 => x"a1c95012",
  1417 => x"c0c4c14a",
  1418 => x"ca501248",
  1419 => x"d8f1c181",
  1420 => x"73501148",
  1421 => x"87f5f849",
  1422 => x"4f264b26",
  1423 => x"c049c01e",
  1424 => x"2687caf7",
  1425 => x"4a711e4f",
  1426 => x"c191cc49",
  1427 => x"c881e0f1",
  1428 => x"c8f4c281",
  1429 => x"c0501148",
  1430 => x"fe49a2f0",
  1431 => x"c087cfed",
  1432 => x"87c3d549",
  1433 => x"ff1e4f26",
  1434 => x"ffc34ad4",
  1435 => x"48d0ff7a",
  1436 => x"de78e1c0",
  1437 => x"487a717a",
  1438 => x"7028b7c8",
  1439 => x"d048717a",
  1440 => x"7a7028b7",
  1441 => x"b7d84871",
  1442 => x"ff7a7028",
  1443 => x"e0c048d0",
  1444 => x"0e4f2678",
  1445 => x"5d5c5b5e",
  1446 => x"7186f40e",
  1447 => x"91cc494d",
  1448 => x"81e0f1c1",
  1449 => x"ca4aa1c8",
  1450 => x"a6c47ea1",
  1451 => x"c4f4c248",
  1452 => x"976e78bf",
  1453 => x"66c44bbf",
  1454 => x"122c734c",
  1455 => x"58a6cc48",
  1456 => x"84c19c70",
  1457 => x"699781c9",
  1458 => x"04acb749",
  1459 => x"4cc087c2",
  1460 => x"4abf976e",
  1461 => x"724966c8",
  1462 => x"c4b9ff31",
  1463 => x"48749966",
  1464 => x"4a703072",
  1465 => x"c8f4c2b1",
  1466 => x"f9fd7159",
  1467 => x"c21ec787",
  1468 => x"1ebfd8f5",
  1469 => x"1ee0f1c1",
  1470 => x"97c8f4c2",
  1471 => x"f4c149bf",
  1472 => x"c0497587",
  1473 => x"e887e5f2",
  1474 => x"264d268e",
  1475 => x"264b264c",
  1476 => x"1e731e4f",
  1477 => x"fd494b71",
  1478 => x"497387f9",
  1479 => x"2687f4fd",
  1480 => x"1e4f264b",
  1481 => x"4b711e73",
  1482 => x"024aa3c2",
  1483 => x"8ac187d6",
  1484 => x"87e2c005",
  1485 => x"bfd8f5c2",
  1486 => x"4887db02",
  1487 => x"f5c288c1",
  1488 => x"87d258dc",
  1489 => x"bfdcf5c2",
  1490 => x"c287cb02",
  1491 => x"48bfd8f5",
  1492 => x"f5c280c1",
  1493 => x"1ec758dc",
  1494 => x"bfd8f5c2",
  1495 => x"e0f1c11e",
  1496 => x"c8f4c21e",
  1497 => x"cc49bf97",
  1498 => x"c0497387",
  1499 => x"f487fdf0",
  1500 => x"264b268e",
  1501 => x"5b5e0e4f",
  1502 => x"ff0e5d5c",
  1503 => x"e8c086cc",
  1504 => x"a6cc59a6",
  1505 => x"c478c048",
  1506 => x"c478c080",
  1507 => x"c478c080",
  1508 => x"66c8c180",
  1509 => x"c180c478",
  1510 => x"c180c478",
  1511 => x"dcf5c278",
  1512 => x"ff78c148",
  1513 => x"e087f6df",
  1514 => x"dfff87d0",
  1515 => x"4d7087e6",
  1516 => x"02adfbc0",
  1517 => x"c087f3c1",
  1518 => x"c10566e4",
  1519 => x"c4c187e8",
  1520 => x"82c44a66",
  1521 => x"cac17e6a",
  1522 => x"496e48dc",
  1523 => x"41204120",
  1524 => x"c4c15110",
  1525 => x"d8c14866",
  1526 => x"496a78cd",
  1527 => x"517581c7",
  1528 => x"4966c4c1",
  1529 => x"51c181c8",
  1530 => x"c248a6dc",
  1531 => x"66c4c178",
  1532 => x"c081c949",
  1533 => x"66c4c151",
  1534 => x"c081ca49",
  1535 => x"d81ec151",
  1536 => x"c8496a1e",
  1537 => x"c5dfff81",
  1538 => x"c186c887",
  1539 => x"c04866c8",
  1540 => x"87c701a8",
  1541 => x"c148a6d4",
  1542 => x"c187cf78",
  1543 => x"c14866c8",
  1544 => x"58a6dc88",
  1545 => x"deff87c4",
  1546 => x"9d7587d0",
  1547 => x"87f1cb02",
  1548 => x"c14866d4",
  1549 => x"03a866cc",
  1550 => x"c087e6cb",
  1551 => x"d3ddff7e",
  1552 => x"484d7087",
  1553 => x"c888c6c1",
  1554 => x"987058a6",
  1555 => x"87d6c102",
  1556 => x"c888c948",
  1557 => x"987058a6",
  1558 => x"87d7c502",
  1559 => x"c888c148",
  1560 => x"987058a6",
  1561 => x"87f8c202",
  1562 => x"c888c348",
  1563 => x"987058a6",
  1564 => x"4887cf02",
  1565 => x"a6c888c1",
  1566 => x"02987058",
  1567 => x"c987f4c4",
  1568 => x"f0c087fe",
  1569 => x"cbdcff7e",
  1570 => x"c04d7087",
  1571 => x"c202adec",
  1572 => x"c07e7587",
  1573 => x"cd02adec",
  1574 => x"f7dbff87",
  1575 => x"c04d7087",
  1576 => x"ff05adec",
  1577 => x"e4c087f3",
  1578 => x"eac10566",
  1579 => x"adecc087",
  1580 => x"ff87c402",
  1581 => x"c087dddb",
  1582 => x"dc1eca1e",
  1583 => x"93cc4b66",
  1584 => x"8366ccc1",
  1585 => x"6c4ca3c4",
  1586 => x"c1dcff49",
  1587 => x"de1ec187",
  1588 => x"ff496c1e",
  1589 => x"d087f7db",
  1590 => x"cdd8c186",
  1591 => x"49a3c87b",
  1592 => x"c95166dc",
  1593 => x"e0c049a3",
  1594 => x"a3ca5166",
  1595 => x"dc516e49",
  1596 => x"80c14866",
  1597 => x"58a6e0c0",
  1598 => x"d84866d4",
  1599 => x"cb04a866",
  1600 => x"4866d487",
  1601 => x"a6d880c1",
  1602 => x"87fac758",
  1603 => x"c14866d8",
  1604 => x"58a6dc88",
  1605 => x"ff87efc7",
  1606 => x"7087dfda",
  1607 => x"87e6c74d",
  1608 => x"87d5dcff",
  1609 => x"d058a6d0",
  1610 => x"c606a866",
  1611 => x"48a6d087",
  1612 => x"ff7866cc",
  1613 => x"c087c2dc",
  1614 => x"c105a8ec",
  1615 => x"e4c087f5",
  1616 => x"e5c10566",
  1617 => x"4966d487",
  1618 => x"c4c191cc",
  1619 => x"a1c48166",
  1620 => x"c84c6a4a",
  1621 => x"66cc4aa1",
  1622 => x"c5d9c152",
  1623 => x"f3d8ff79",
  1624 => x"9d4d7087",
  1625 => x"c087da02",
  1626 => x"d402adfb",
  1627 => x"ff547587",
  1628 => x"7087e1d8",
  1629 => x"c0029d4d",
  1630 => x"fbc087c7",
  1631 => x"ecff05ad",
  1632 => x"54e0c087",
  1633 => x"c054c1c2",
  1634 => x"66d47c97",
  1635 => x"a866d848",
  1636 => x"87cbc004",
  1637 => x"c14866d4",
  1638 => x"58a6d880",
  1639 => x"d887e7c5",
  1640 => x"88c14866",
  1641 => x"c558a6dc",
  1642 => x"d8ff87dc",
  1643 => x"4d7087cc",
  1644 => x"cc87d3c5",
  1645 => x"e4c04866",
  1646 => x"c405a866",
  1647 => x"e8c087f4",
  1648 => x"78c048a6",
  1649 => x"87f1d9ff",
  1650 => x"d9ff7e70",
  1651 => x"f0c087eb",
  1652 => x"ecc058a6",
  1653 => x"c7c005a8",
  1654 => x"6e48a687",
  1655 => x"87c4c078",
  1656 => x"87f0d6ff",
  1657 => x"cc4966d4",
  1658 => x"66c4c191",
  1659 => x"c8807148",
  1660 => x"66c458a6",
  1661 => x"c482c84a",
  1662 => x"81ca4966",
  1663 => x"ecc0516e",
  1664 => x"81c14966",
  1665 => x"48c1896e",
  1666 => x"49703071",
  1667 => x"977189c1",
  1668 => x"c4f4c27a",
  1669 => x"296e49bf",
  1670 => x"484a6a97",
  1671 => x"f4c09871",
  1672 => x"66c458a6",
  1673 => x"cc80c448",
  1674 => x"66c858a6",
  1675 => x"e4c04cbf",
  1676 => x"66cc4866",
  1677 => x"c5c002a8",
  1678 => x"c07ec087",
  1679 => x"7ec187c2",
  1680 => x"e0c01e6e",
  1681 => x"ff49741e",
  1682 => x"c887c3d6",
  1683 => x"c04d7086",
  1684 => x"c106adb7",
  1685 => x"847587d4",
  1686 => x"49bf66c8",
  1687 => x"7481e0c0",
  1688 => x"cac14b89",
  1689 => x"fe714ae8",
  1690 => x"c287f7de",
  1691 => x"c07e7484",
  1692 => x"c14866e8",
  1693 => x"a6ecc080",
  1694 => x"66f0c058",
  1695 => x"7081c149",
  1696 => x"c5c002a9",
  1697 => x"c04cc087",
  1698 => x"4cc187c2",
  1699 => x"66cc1e74",
  1700 => x"e0c049bf",
  1701 => x"8966c481",
  1702 => x"66c81e71",
  1703 => x"edd4ff49",
  1704 => x"c086c887",
  1705 => x"ff01a8b7",
  1706 => x"e8c087c5",
  1707 => x"d3c00266",
  1708 => x"4966c487",
  1709 => x"e8c081c9",
  1710 => x"66c45166",
  1711 => x"d3dac148",
  1712 => x"87cec078",
  1713 => x"c94966c4",
  1714 => x"c451c281",
  1715 => x"dcc14866",
  1716 => x"66d478d1",
  1717 => x"a866d848",
  1718 => x"87cbc004",
  1719 => x"c14866d4",
  1720 => x"58a6d880",
  1721 => x"d887d1c0",
  1722 => x"88c14866",
  1723 => x"c058a6dc",
  1724 => x"d3ff87c6",
  1725 => x"4d7087c4",
  1726 => x"c048a6cc",
  1727 => x"87c6c078",
  1728 => x"87f6d2ff",
  1729 => x"e0c04d70",
  1730 => x"80c14866",
  1731 => x"58a6e4c0",
  1732 => x"c0029d75",
  1733 => x"66d487cb",
  1734 => x"66ccc148",
  1735 => x"daf404a8",
  1736 => x"4866d487",
  1737 => x"c003a8c7",
  1738 => x"66d487e1",
  1739 => x"dcf5c24c",
  1740 => x"7478c048",
  1741 => x"c191cc49",
  1742 => x"c48166c4",
  1743 => x"4a6a4aa1",
  1744 => x"c17952c0",
  1745 => x"04acc784",
  1746 => x"c087e2ff",
  1747 => x"c00266e4",
  1748 => x"c4c187e2",
  1749 => x"d4c14966",
  1750 => x"66c4c181",
  1751 => x"82dcc14a",
  1752 => x"d9c152c0",
  1753 => x"c4c179c5",
  1754 => x"d8c14966",
  1755 => x"eccac181",
  1756 => x"87d6c079",
  1757 => x"4966c4c1",
  1758 => x"c181d4c1",
  1759 => x"c14a66c4",
  1760 => x"cac182d8",
  1761 => x"d8c17af4",
  1762 => x"c4c179fc",
  1763 => x"e0c14966",
  1764 => x"e3dcc181",
  1765 => x"d8d0ff79",
  1766 => x"4866d087",
  1767 => x"268eccff",
  1768 => x"264c264d",
  1769 => x"1e4f264b",
  1770 => x"f5c21ec7",
  1771 => x"c11ebfd8",
  1772 => x"c21ee0f1",
  1773 => x"bf97c8f4",
  1774 => x"87f9ee49",
  1775 => x"49e0f1c1",
  1776 => x"87f6e0c0",
  1777 => x"4f268ef4",
  1778 => x"d4f1c11e",
  1779 => x"c150c048",
  1780 => x"49bfccf3",
  1781 => x"87ced5ff",
  1782 => x"4f2648c0",
  1783 => x"c71e731e",
  1784 => x"f5c287cc",
  1785 => x"50c048e4",
  1786 => x"c348d4ff",
  1787 => x"cac178ff",
  1788 => x"d7fe49fc",
  1789 => x"e2fe87d3",
  1790 => x"987087e6",
  1791 => x"fe87cd02",
  1792 => x"7087c4ec",
  1793 => x"87c40298",
  1794 => x"87c24ac1",
  1795 => x"9a724ac0",
  1796 => x"c187c802",
  1797 => x"fe49c8cb",
  1798 => x"c287eed6",
  1799 => x"c048d8f5",
  1800 => x"c8f4c278",
  1801 => x"4950c048",
  1802 => x"fe87fcfd",
  1803 => x"4b7087da",
  1804 => x"87ce029b",
  1805 => x"5bfcf2c1",
  1806 => x"efdd49c7",
  1807 => x"df49c187",
  1808 => x"f2c287cb",
  1809 => x"d1e0c087",
  1810 => x"e3eec087",
  1811 => x"87f5ff87",
  1812 => x"4f264b26",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"00000001",
  1816 => x"0000131e",
  1817 => x"00002d70",
  1818 => x"54000000",
  1819 => x"0000131e",
  1820 => x"00002d8e",
  1821 => x"54000000",
  1822 => x"0000131e",
  1823 => x"00002dac",
  1824 => x"54000000",
  1825 => x"0000131e",
  1826 => x"00002dca",
  1827 => x"54000000",
  1828 => x"0000131e",
  1829 => x"00002de8",
  1830 => x"54000000",
  1831 => x"0000131e",
  1832 => x"00002e06",
  1833 => x"54000000",
  1834 => x"0000131e",
  1835 => x"00002e24",
  1836 => x"54000000",
  1837 => x"00001645",
  1838 => x"00000000",
  1839 => x"54000000",
  1840 => x"000013f7",
  1841 => x"00000000",
  1842 => x"54000000",
  1843 => x"000012cc",
  1844 => x"db86fc1e",
  1845 => x"fc7e7087",
  1846 => x"1e4f268e",
  1847 => x"c048f0fe",
  1848 => x"7909cd78",
  1849 => x"1e4f2609",
  1850 => x"49d0f3c1",
  1851 => x"4f2687ed",
  1852 => x"bff0fe1e",
  1853 => x"1e4f2648",
  1854 => x"c148f0fe",
  1855 => x"1e4f2678",
  1856 => x"c048f0fe",
  1857 => x"1e4f2678",
  1858 => x"52c04a71",
  1859 => x"0e4f2651",
  1860 => x"5d5c5b5e",
  1861 => x"7186f40e",
  1862 => x"7e6d974d",
  1863 => x"974ca5c1",
  1864 => x"a6c8486c",
  1865 => x"c4486e58",
  1866 => x"c505a866",
  1867 => x"c048ff87",
  1868 => x"caff87e6",
  1869 => x"49a5c287",
  1870 => x"714b6c97",
  1871 => x"6b974ba3",
  1872 => x"7e6c974b",
  1873 => x"80c1486e",
  1874 => x"c758a6c8",
  1875 => x"58a6cc98",
  1876 => x"fe7c9770",
  1877 => x"487387e1",
  1878 => x"4d268ef4",
  1879 => x"4b264c26",
  1880 => x"731e4f26",
  1881 => x"fe86f41e",
  1882 => x"bfe087d5",
  1883 => x"e0c0494b",
  1884 => x"c00299c0",
  1885 => x"4a7387ea",
  1886 => x"c29affc3",
  1887 => x"bf97d8f9",
  1888 => x"daf9c249",
  1889 => x"c2517281",
  1890 => x"bf97d8f9",
  1891 => x"c1486e7e",
  1892 => x"58a6c880",
  1893 => x"a6cc98c7",
  1894 => x"d8f9c258",
  1895 => x"5066c848",
  1896 => x"7087cdfd",
  1897 => x"87cffd7e",
  1898 => x"4b268ef4",
  1899 => x"c21e4f26",
  1900 => x"fd49d8f9",
  1901 => x"f5c187d1",
  1902 => x"defc49e2",
  1903 => x"87f0c387",
  1904 => x"731e4f26",
  1905 => x"d8f9c21e",
  1906 => x"87c3fd49",
  1907 => x"b7c04a70",
  1908 => x"ccc204aa",
  1909 => x"aaf0c387",
  1910 => x"c187c905",
  1911 => x"c148e8f9",
  1912 => x"87edc178",
  1913 => x"05aae0c3",
  1914 => x"f9c187c9",
  1915 => x"78c148ec",
  1916 => x"c187dec1",
  1917 => x"02bfecf9",
  1918 => x"c0c287c6",
  1919 => x"87c24ba2",
  1920 => x"f9c14b72",
  1921 => x"c002bfe8",
  1922 => x"497387e0",
  1923 => x"9129b7c4",
  1924 => x"81f0f9c1",
  1925 => x"9acf4a73",
  1926 => x"48c192c2",
  1927 => x"4a703072",
  1928 => x"4872baff",
  1929 => x"79709869",
  1930 => x"497387db",
  1931 => x"9129b7c4",
  1932 => x"81f0f9c1",
  1933 => x"9acf4a73",
  1934 => x"48c392c2",
  1935 => x"4a703072",
  1936 => x"70b06948",
  1937 => x"ecf9c179",
  1938 => x"c178c048",
  1939 => x"c048e8f9",
  1940 => x"d8f9c278",
  1941 => x"87f7fa49",
  1942 => x"b7c04a70",
  1943 => x"f4fd03aa",
  1944 => x"2648c087",
  1945 => x"004f264b",
  1946 => x"00000000",
  1947 => x"00000000",
  1948 => x"00000000",
  1949 => x"84848484",
  1950 => x"84848484",
  1951 => x"84848484",
  1952 => x"84848484",
  1953 => x"84848484",
  1954 => x"84848484",
  1955 => x"84848484",
  1956 => x"84848484",
  1957 => x"84848484",
  1958 => x"84848484",
  1959 => x"84848484",
  1960 => x"84848484",
  1961 => x"84848484",
  1962 => x"84848484",
  1963 => x"84848484",
  1964 => x"724ac01e",
  1965 => x"c191c449",
  1966 => x"c081f0f9",
  1967 => x"d082c179",
  1968 => x"ee04aab7",
  1969 => x"0e4f2687",
  1970 => x"5d5c5b5e",
  1971 => x"f84d710e",
  1972 => x"4a7587ed",
  1973 => x"922ab7c4",
  1974 => x"82f0f9c1",
  1975 => x"9ccf4c75",
  1976 => x"496a94c2",
  1977 => x"c32b744b",
  1978 => x"7448c29b",
  1979 => x"ff4c7030",
  1980 => x"714874bc",
  1981 => x"f77a7098",
  1982 => x"487387fd",
  1983 => x"4c264d26",
  1984 => x"4f264b26",
  1985 => x"48d0ff1e",
  1986 => x"7178e1c8",
  1987 => x"08d4ff48",
  1988 => x"1e4f2678",
  1989 => x"c848d0ff",
  1990 => x"487178e1",
  1991 => x"7808d4ff",
  1992 => x"ff4866c4",
  1993 => x"267808d4",
  1994 => x"4a711e4f",
  1995 => x"1e4966c4",
  1996 => x"deff4972",
  1997 => x"48d0ff87",
  1998 => x"fc78e0c0",
  1999 => x"1e4f268e",
  2000 => x"4b711e73",
  2001 => x"1e4966c8",
  2002 => x"e0c14a73",
  2003 => x"d8ff49a2",
  2004 => x"268efc87",
  2005 => x"1e4f264b",
  2006 => x"c848d0ff",
  2007 => x"487178c9",
  2008 => x"7808d4ff",
  2009 => x"711e4f26",
  2010 => x"87eb494a",
  2011 => x"c848d0ff",
  2012 => x"1e4f2678",
  2013 => x"4b711e73",
  2014 => x"bff0f9c2",
  2015 => x"c287c302",
  2016 => x"d0ff87eb",
  2017 => x"78c9c848",
  2018 => x"e0c04873",
  2019 => x"08d4ffb0",
  2020 => x"e4f9c278",
  2021 => x"c878c048",
  2022 => x"87c50266",
  2023 => x"c249ffc3",
  2024 => x"c249c087",
  2025 => x"cc59ecf9",
  2026 => x"87c60266",
  2027 => x"4ad5d5c5",
  2028 => x"ffcf87c4",
  2029 => x"f9c24aff",
  2030 => x"f9c25af0",
  2031 => x"78c148f0",
  2032 => x"4f264b26",
  2033 => x"5c5b5e0e",
  2034 => x"4d710e5d",
  2035 => x"bfecf9c2",
  2036 => x"029d754b",
  2037 => x"c84987cb",
  2038 => x"ecfdc191",
  2039 => x"c482714a",
  2040 => x"ecc1c287",
  2041 => x"124cc04a",
  2042 => x"c2997349",
  2043 => x"48bfe8f9",
  2044 => x"d4ffb871",
  2045 => x"b7c17808",
  2046 => x"b7c8842b",
  2047 => x"87e704ac",
  2048 => x"bfe4f9c2",
  2049 => x"c280c848",
  2050 => x"2658e8f9",
  2051 => x"264c264d",
  2052 => x"1e4f264b",
  2053 => x"4b711e73",
  2054 => x"029a4a13",
  2055 => x"497287cb",
  2056 => x"1387e1fe",
  2057 => x"f5059a4a",
  2058 => x"264b2687",
  2059 => x"f9c21e4f",
  2060 => x"c249bfe4",
  2061 => x"c148e4f9",
  2062 => x"c0c478a1",
  2063 => x"db03a9b7",
  2064 => x"48d4ff87",
  2065 => x"bfe8f9c2",
  2066 => x"e4f9c278",
  2067 => x"f9c249bf",
  2068 => x"a1c148e4",
  2069 => x"b7c0c478",
  2070 => x"87e504a9",
  2071 => x"c848d0ff",
  2072 => x"f0f9c278",
  2073 => x"2678c048",
  2074 => x"0000004f",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"5f000000",
  2078 => x"0000005f",
  2079 => x"00030300",
  2080 => x"00000303",
  2081 => x"147f7f14",
  2082 => x"00147f7f",
  2083 => x"6b2e2400",
  2084 => x"00123a6b",
  2085 => x"18366a4c",
  2086 => x"0032566c",
  2087 => x"594f7e30",
  2088 => x"40683a77",
  2089 => x"07040000",
  2090 => x"00000003",
  2091 => x"3e1c0000",
  2092 => x"00004163",
  2093 => x"63410000",
  2094 => x"00001c3e",
  2095 => x"1c3e2a08",
  2096 => x"082a3e1c",
  2097 => x"3e080800",
  2098 => x"0008083e",
  2099 => x"e0800000",
  2100 => x"00000060",
  2101 => x"08080800",
  2102 => x"00080808",
  2103 => x"60000000",
  2104 => x"00000060",
  2105 => x"18306040",
  2106 => x"0103060c",
  2107 => x"597f3e00",
  2108 => x"003e7f4d",
  2109 => x"7f060400",
  2110 => x"0000007f",
  2111 => x"71634200",
  2112 => x"00464f59",
  2113 => x"49632200",
  2114 => x"00367f49",
  2115 => x"13161c18",
  2116 => x"00107f7f",
  2117 => x"45672700",
  2118 => x"00397d45",
  2119 => x"4b7e3c00",
  2120 => x"00307949",
  2121 => x"71010100",
  2122 => x"00070f79",
  2123 => x"497f3600",
  2124 => x"00367f49",
  2125 => x"494f0600",
  2126 => x"001e3f69",
  2127 => x"66000000",
  2128 => x"00000066",
  2129 => x"e6800000",
  2130 => x"00000066",
  2131 => x"14080800",
  2132 => x"00222214",
  2133 => x"14141400",
  2134 => x"00141414",
  2135 => x"14222200",
  2136 => x"00080814",
  2137 => x"51030200",
  2138 => x"00060f59",
  2139 => x"5d417f3e",
  2140 => x"001e1f55",
  2141 => x"097f7e00",
  2142 => x"007e7f09",
  2143 => x"497f7f00",
  2144 => x"00367f49",
  2145 => x"633e1c00",
  2146 => x"00414141",
  2147 => x"417f7f00",
  2148 => x"001c3e63",
  2149 => x"497f7f00",
  2150 => x"00414149",
  2151 => x"097f7f00",
  2152 => x"00010109",
  2153 => x"417f3e00",
  2154 => x"007a7b49",
  2155 => x"087f7f00",
  2156 => x"007f7f08",
  2157 => x"7f410000",
  2158 => x"0000417f",
  2159 => x"40602000",
  2160 => x"003f7f40",
  2161 => x"1c087f7f",
  2162 => x"00416336",
  2163 => x"407f7f00",
  2164 => x"00404040",
  2165 => x"0c067f7f",
  2166 => x"007f7f06",
  2167 => x"0c067f7f",
  2168 => x"007f7f18",
  2169 => x"417f3e00",
  2170 => x"003e7f41",
  2171 => x"097f7f00",
  2172 => x"00060f09",
  2173 => x"61417f3e",
  2174 => x"00407e7f",
  2175 => x"097f7f00",
  2176 => x"00667f19",
  2177 => x"4d6f2600",
  2178 => x"00327b59",
  2179 => x"7f010100",
  2180 => x"0001017f",
  2181 => x"407f3f00",
  2182 => x"003f7f40",
  2183 => x"703f0f00",
  2184 => x"000f3f70",
  2185 => x"18307f7f",
  2186 => x"007f7f30",
  2187 => x"1c366341",
  2188 => x"4163361c",
  2189 => x"7c060301",
  2190 => x"0103067c",
  2191 => x"4d597161",
  2192 => x"00414347",
  2193 => x"7f7f0000",
  2194 => x"00004141",
  2195 => x"0c060301",
  2196 => x"40603018",
  2197 => x"41410000",
  2198 => x"00007f7f",
  2199 => x"03060c08",
  2200 => x"00080c06",
  2201 => x"80808080",
  2202 => x"00808080",
  2203 => x"03000000",
  2204 => x"00000407",
  2205 => x"54742000",
  2206 => x"00787c54",
  2207 => x"447f7f00",
  2208 => x"00387c44",
  2209 => x"447c3800",
  2210 => x"00004444",
  2211 => x"447c3800",
  2212 => x"007f7f44",
  2213 => x"547c3800",
  2214 => x"00185c54",
  2215 => x"7f7e0400",
  2216 => x"00000505",
  2217 => x"a4bc1800",
  2218 => x"007cfca4",
  2219 => x"047f7f00",
  2220 => x"00787c04",
  2221 => x"3d000000",
  2222 => x"0000407d",
  2223 => x"80808000",
  2224 => x"00007dfd",
  2225 => x"107f7f00",
  2226 => x"00446c38",
  2227 => x"3f000000",
  2228 => x"0000407f",
  2229 => x"180c7c7c",
  2230 => x"00787c0c",
  2231 => x"047c7c00",
  2232 => x"00787c04",
  2233 => x"447c3800",
  2234 => x"00387c44",
  2235 => x"24fcfc00",
  2236 => x"00183c24",
  2237 => x"243c1800",
  2238 => x"00fcfc24",
  2239 => x"047c7c00",
  2240 => x"00080c04",
  2241 => x"545c4800",
  2242 => x"00207454",
  2243 => x"7f3f0400",
  2244 => x"00004444",
  2245 => x"407c3c00",
  2246 => x"007c7c40",
  2247 => x"603c1c00",
  2248 => x"001c3c60",
  2249 => x"30607c3c",
  2250 => x"003c7c60",
  2251 => x"10386c44",
  2252 => x"00446c38",
  2253 => x"e0bc1c00",
  2254 => x"001c3c60",
  2255 => x"74644400",
  2256 => x"00444c5c",
  2257 => x"3e080800",
  2258 => x"00414177",
  2259 => x"7f000000",
  2260 => x"0000007f",
  2261 => x"77414100",
  2262 => x"0008083e",
  2263 => x"03010102",
  2264 => x"00010202",
  2265 => x"7f7f7f7f",
  2266 => x"007f7f7f",
  2267 => x"1c1c0808",
  2268 => x"7f7f3e3e",
  2269 => x"3e3e7f7f",
  2270 => x"08081c1c",
  2271 => x"7c181000",
  2272 => x"0010187c",
  2273 => x"7c301000",
  2274 => x"0010307c",
  2275 => x"60603010",
  2276 => x"00061e78",
  2277 => x"183c6642",
  2278 => x"0042663c",
  2279 => x"c26a3878",
  2280 => x"00386cc6",
  2281 => x"60000060",
  2282 => x"00600000",
  2283 => x"5c5b5e0e",
  2284 => x"86fc0e5d",
  2285 => x"f9c27e71",
  2286 => x"c04cbff8",
  2287 => x"c41ec04b",
  2288 => x"c402ab66",
  2289 => x"c24dc087",
  2290 => x"754dc187",
  2291 => x"ee49731e",
  2292 => x"86c887e1",
  2293 => x"ef49e0c0",
  2294 => x"a4c487ea",
  2295 => x"f0496a4a",
  2296 => x"c8f187f1",
  2297 => x"c184cc87",
  2298 => x"abb7c883",
  2299 => x"87cdff04",
  2300 => x"4d268efc",
  2301 => x"4b264c26",
  2302 => x"711e4f26",
  2303 => x"fcf9c24a",
  2304 => x"fcf9c25a",
  2305 => x"4978c748",
  2306 => x"2687e1fe",
  2307 => x"1e731e4f",
  2308 => x"0bfc4b71",
  2309 => x"4a730b7b",
  2310 => x"c0c19ac1",
  2311 => x"c5ed49a2",
  2312 => x"fcddc287",
  2313 => x"264b265b",
  2314 => x"4a711e4f",
  2315 => x"721e66c4",
  2316 => x"87cbec49",
  2317 => x"4f268efc",
  2318 => x"48d4ff1e",
  2319 => x"ff78ffc3",
  2320 => x"e1c048d0",
  2321 => x"48d4ff78",
  2322 => x"487178c1",
  2323 => x"d4ff30c4",
  2324 => x"d0ff7808",
  2325 => x"78e0c048",
  2326 => x"5e0e4f26",
  2327 => x"0e5d5c5b",
  2328 => x"a6c886ec",
  2329 => x"c478c048",
  2330 => x"78bfec80",
  2331 => x"f9c280f8",
  2332 => x"c278bff8",
  2333 => x"4cbfc0fa",
  2334 => x"c24dbfe8",
  2335 => x"49bff8dd",
  2336 => x"c787ffe4",
  2337 => x"87ffe849",
  2338 => x"99c24970",
  2339 => x"c287d005",
  2340 => x"49bff0dd",
  2341 => x"66ccb9ff",
  2342 => x"0299c199",
  2343 => x"c887cbc2",
  2344 => x"c8ff48a6",
  2345 => x"49c778bf",
  2346 => x"7087dce8",
  2347 => x"717e7449",
  2348 => x"87cd0599",
  2349 => x"c14966cc",
  2350 => x"717e7499",
  2351 => x"c4c10299",
  2352 => x"4cc8ff87",
  2353 => x"cc4b66c8",
  2354 => x"bfec48a6",
  2355 => x"87f2e378",
  2356 => x"6c5ba6cc",
  2357 => x"d4887348",
  2358 => x"e8cf58a6",
  2359 => x"87d106a8",
  2360 => x"bfecddc2",
  2361 => x"c2b9c149",
  2362 => x"7159f0dd",
  2363 => x"6c87c9fd",
  2364 => x"e749c74b",
  2365 => x"987087d1",
  2366 => x"87cbff05",
  2367 => x"c14966cc",
  2368 => x"c2ff0599",
  2369 => x"c24c6e87",
  2370 => x"4abff8dd",
  2371 => x"ddc2bac1",
  2372 => x"0afc5afc",
  2373 => x"9ac10a7a",
  2374 => x"49a2c0c1",
  2375 => x"c187c7e9",
  2376 => x"e2e649da",
  2377 => x"48a6c887",
  2378 => x"ddc278c1",
  2379 => x"66cc48f0",
  2380 => x"f8ddc278",
  2381 => x"c7c105bf",
  2382 => x"c0c0c887",
  2383 => x"dcddc24b",
  2384 => x"144c6e7e",
  2385 => x"87ffe549",
  2386 => x"c0029870",
  2387 => x"b57387c2",
  2388 => x"052bb7c1",
  2389 => x"7587ecff",
  2390 => x"99ffc349",
  2391 => x"49c01e71",
  2392 => x"7587c6fb",
  2393 => x"29b7c849",
  2394 => x"49c11e71",
  2395 => x"c887fafa",
  2396 => x"49fdc386",
  2397 => x"c387d0e5",
  2398 => x"cae549fa",
  2399 => x"87cec787",
  2400 => x"ffc34975",
  2401 => x"2db7c899",
  2402 => x"9d75b571",
  2403 => x"87e0c002",
  2404 => x"7ebfc8ff",
  2405 => x"ddc2496e",
  2406 => x"c289bff4",
  2407 => x"c003a9e0",
  2408 => x"4dc087c5",
  2409 => x"c287cfc0",
  2410 => x"6e48f4dd",
  2411 => x"87c6c078",
  2412 => x"48f4ddc2",
  2413 => x"497578c0",
  2414 => x"c00599c8",
  2415 => x"f5c387ce",
  2416 => x"87c3e449",
  2417 => x"99c24970",
  2418 => x"87eac002",
  2419 => x"bffcf9c2",
  2420 => x"87cac002",
  2421 => x"c288c148",
  2422 => x"c058c0fa",
  2423 => x"66c487d3",
  2424 => x"80e0c148",
  2425 => x"bf6e7e70",
  2426 => x"87c5c002",
  2427 => x"7349ff4b",
  2428 => x"48a6c80f",
  2429 => x"497578c1",
  2430 => x"c00599c4",
  2431 => x"f2c387ce",
  2432 => x"87c3e349",
  2433 => x"99c24970",
  2434 => x"87f1c002",
  2435 => x"bffcf9c2",
  2436 => x"c7486e7e",
  2437 => x"c003a8b7",
  2438 => x"486e87cb",
  2439 => x"fac280c1",
  2440 => x"d3c058c0",
  2441 => x"4866c487",
  2442 => x"7080e0c1",
  2443 => x"02bf6e7e",
  2444 => x"4b87c5c0",
  2445 => x"0f7349fe",
  2446 => x"c148a6c8",
  2447 => x"49fdc378",
  2448 => x"7087c4e2",
  2449 => x"0299c249",
  2450 => x"c287e6c0",
  2451 => x"02bffcf9",
  2452 => x"c287c9c0",
  2453 => x"c048fcf9",
  2454 => x"87d0c078",
  2455 => x"c14a66c4",
  2456 => x"026a82e0",
  2457 => x"4b87c5c0",
  2458 => x"0f7349fd",
  2459 => x"c148a6c8",
  2460 => x"49fac378",
  2461 => x"7087d0e1",
  2462 => x"0299c249",
  2463 => x"c287edc0",
  2464 => x"48bffcf9",
  2465 => x"03a8b7c7",
  2466 => x"c287c9c0",
  2467 => x"c748fcf9",
  2468 => x"87d3c078",
  2469 => x"c14866c4",
  2470 => x"7e7080e0",
  2471 => x"c002bf6e",
  2472 => x"fc4b87c5",
  2473 => x"c80f7349",
  2474 => x"78c148a6",
  2475 => x"f0c34875",
  2476 => x"487e7098",
  2477 => x"cec00598",
  2478 => x"49dac187",
  2479 => x"7087c8e0",
  2480 => x"0299c249",
  2481 => x"6e87cac1",
  2482 => x"87cdc005",
  2483 => x"ff49dac1",
  2484 => x"7087f4df",
  2485 => x"e8c00298",
  2486 => x"49bfe887",
  2487 => x"9bffc34b",
  2488 => x"7129b7c8",
  2489 => x"d9dbffb3",
  2490 => x"c3497387",
  2491 => x"997199f0",
  2492 => x"87e5ff05",
  2493 => x"ff49dac1",
  2494 => x"7087ccdf",
  2495 => x"d8ff0598",
  2496 => x"fcf9c287",
  2497 => x"cc4b49bf",
  2498 => x"8366c493",
  2499 => x"73714b6b",
  2500 => x"029c740f",
  2501 => x"6c87e9c0",
  2502 => x"87e4c002",
  2503 => x"deff496c",
  2504 => x"497087e5",
  2505 => x"c00299c1",
  2506 => x"a4c487cb",
  2507 => x"fcf9c24b",
  2508 => x"4b6b49bf",
  2509 => x"0284c80f",
  2510 => x"6c87c5c0",
  2511 => x"87dcff05",
  2512 => x"c00266c8",
  2513 => x"f9c287c8",
  2514 => x"f149bffc",
  2515 => x"8eec87de",
  2516 => x"4c264d26",
  2517 => x"4f264b26",
  2518 => x"00000010",
  2519 => x"14111258",
  2520 => x"231c1b1d",
  2521 => x"9491595a",
  2522 => x"f4ebf2f5",
  2523 => x"00000000",
  2524 => x"00000000",
  2525 => x"00000000",
  2526 => x"00000000",
  2527 => x"5c5b5e0e",
  2528 => x"4b710e5d",
  2529 => x"d04cd4ff",
  2530 => x"78c04866",
  2531 => x"ddff49d6",
  2532 => x"ffc387f2",
  2533 => x"c3496c7c",
  2534 => x"4d7199ff",
  2535 => x"99f0c349",
  2536 => x"05a9e0c1",
  2537 => x"ffc387cb",
  2538 => x"c3486c7c",
  2539 => x"0866d098",
  2540 => x"7cffc378",
  2541 => x"c8494a6c",
  2542 => x"7cffc331",
  2543 => x"b2714a6c",
  2544 => x"31c84972",
  2545 => x"6c7cffc3",
  2546 => x"72b2714a",
  2547 => x"c331c849",
  2548 => x"4a6c7cff",
  2549 => x"d0ffb271",
  2550 => x"78e0c048",
  2551 => x"c2029b73",
  2552 => x"757b7287",
  2553 => x"264d2648",
  2554 => x"264b264c",
  2555 => x"4f261e4f",
  2556 => x"5c5b5e0e",
  2557 => x"7686f80e",
  2558 => x"49a6c81e",
  2559 => x"c487fdfd",
  2560 => x"6e4b7086",
  2561 => x"01a8c348",
  2562 => x"7387f4c2",
  2563 => x"9af0c34a",
  2564 => x"02aad0c1",
  2565 => x"e0c187c7",
  2566 => x"e2c205aa",
  2567 => x"c8497387",
  2568 => x"87c30299",
  2569 => x"7387c6ff",
  2570 => x"c29cc34c",
  2571 => x"c4c105ac",
  2572 => x"4966c487",
  2573 => x"1e7131c9",
  2574 => x"c14a66c4",
  2575 => x"fac292cc",
  2576 => x"817249c4",
  2577 => x"87e6cefe",
  2578 => x"daff49d8",
  2579 => x"c0c887f6",
  2580 => x"fce6c21e",
  2581 => x"fce7fd49",
  2582 => x"48d0ff87",
  2583 => x"c278e0c0",
  2584 => x"cc1efce6",
  2585 => x"ccc14a66",
  2586 => x"c4fac292",
  2587 => x"fe817249",
  2588 => x"cc87fccc",
  2589 => x"05acc186",
  2590 => x"c487c4c1",
  2591 => x"31c94966",
  2592 => x"66c41e71",
  2593 => x"92ccc14a",
  2594 => x"49c4fac2",
  2595 => x"cdfe8172",
  2596 => x"e6c287dc",
  2597 => x"66c81efc",
  2598 => x"92ccc14a",
  2599 => x"49c4fac2",
  2600 => x"cbfe8172",
  2601 => x"49d787ca",
  2602 => x"87d8d9ff",
  2603 => x"c21ec0c8",
  2604 => x"fd49fce6",
  2605 => x"cc87fbe5",
  2606 => x"48d0ff86",
  2607 => x"f878e0c0",
  2608 => x"264c268e",
  2609 => x"1e4f264b",
  2610 => x"b7c44a71",
  2611 => x"87ce03aa",
  2612 => x"ccc14972",
  2613 => x"c4fac291",
  2614 => x"81c8c181",
  2615 => x"4f2679c0",
  2616 => x"5c5b5e0e",
  2617 => x"86fc0e5d",
  2618 => x"d4ff4a71",
  2619 => x"d44cc04b",
  2620 => x"b7c34d66",
  2621 => x"c2c201ad",
  2622 => x"029a7287",
  2623 => x"1e87ecc0",
  2624 => x"ccc14975",
  2625 => x"c4fac291",
  2626 => x"c8807148",
  2627 => x"66c458a6",
  2628 => x"e7c4fe49",
  2629 => x"7086c487",
  2630 => x"87d40298",
  2631 => x"c8c1496e",
  2632 => x"6e79c181",
  2633 => x"6981c849",
  2634 => x"7587c54c",
  2635 => x"87d7fe49",
  2636 => x"c848d0ff",
  2637 => x"7bdd78e1",
  2638 => x"ffc34874",
  2639 => x"747b7098",
  2640 => x"29b7c849",
  2641 => x"ffc34871",
  2642 => x"747b7098",
  2643 => x"29b7d049",
  2644 => x"ffc34871",
  2645 => x"747b7098",
  2646 => x"28b7d848",
  2647 => x"7bc07b70",
  2648 => x"7b7b7b7b",
  2649 => x"7b7b7b7b",
  2650 => x"ff7b7b7b",
  2651 => x"e0c048d0",
  2652 => x"dc1e7578",
  2653 => x"f0d6ff49",
  2654 => x"fc86c487",
  2655 => x"264d268e",
  2656 => x"264b264c",
  2657 => x"001ce74f",
  2658 => x"001ce700",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
