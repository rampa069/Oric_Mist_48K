
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"fe",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"f4",x"fe",x"c2"),
    18 => (x"48",x"cc",x"e6",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"c9",x"e6",x"c2",x"87"),
    25 => (x"c5",x"e6",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"ed",x"c1",x"87",x"f7"),
    29 => (x"e6",x"c2",x"87",x"e6"),
    30 => (x"e6",x"c2",x"4d",x"c9"),
    31 => (x"ad",x"74",x"4c",x"c9"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"86",x"f0",x"0e",x"5d"),
    37 => (x"a6",x"c4",x"4c",x"c0"),
    38 => (x"c0",x"78",x"c0",x"48"),
    39 => (x"c0",x"4b",x"a6",x"e4"),
    40 => (x"48",x"49",x"66",x"e0"),
    41 => (x"e4",x"c0",x"80",x"c1"),
    42 => (x"7e",x"11",x"58",x"a6"),
    43 => (x"f1",x"c3",x"02",x"6e"),
    44 => (x"02",x"66",x"c4",x"87"),
    45 => (x"c4",x"87",x"c6",x"c3"),
    46 => (x"78",x"c0",x"48",x"a6"),
    47 => (x"f0",x"c0",x"4a",x"6e"),
    48 => (x"da",x"c2",x"02",x"8a"),
    49 => (x"8a",x"f3",x"c0",x"87"),
    50 => (x"87",x"db",x"c2",x"02"),
    51 => (x"dc",x"02",x"8a",x"c1"),
    52 => (x"02",x"8a",x"c8",x"87"),
    53 => (x"c4",x"87",x"c8",x"c2"),
    54 => (x"87",x"d1",x"02",x"8a"),
    55 => (x"c1",x"02",x"8a",x"c3"),
    56 => (x"8a",x"c2",x"87",x"eb"),
    57 => (x"c3",x"87",x"c6",x"02"),
    58 => (x"c9",x"c2",x"05",x"8a"),
    59 => (x"73",x"83",x"c4",x"87"),
    60 => (x"69",x"89",x"c4",x"49"),
    61 => (x"c1",x"02",x"6e",x"7e"),
    62 => (x"a6",x"c8",x"87",x"c8"),
    63 => (x"c4",x"78",x"c0",x"48"),
    64 => (x"cc",x"78",x"c0",x"80"),
    65 => (x"4a",x"6e",x"4d",x"66"),
    66 => (x"cf",x"2a",x"b7",x"dc"),
    67 => (x"c4",x"48",x"6e",x"9a"),
    68 => (x"72",x"7e",x"70",x"30"),
    69 => (x"87",x"c5",x"02",x"9a"),
    70 => (x"c1",x"48",x"a6",x"c8"),
    71 => (x"06",x"aa",x"c9",x"78"),
    72 => (x"f7",x"c0",x"87",x"c5"),
    73 => (x"c0",x"87",x"c3",x"82"),
    74 => (x"66",x"c8",x"82",x"f0"),
    75 => (x"72",x"87",x"c7",x"02"),
    76 => (x"87",x"fa",x"c1",x"49"),
    77 => (x"85",x"c1",x"84",x"c1"),
    78 => (x"04",x"ad",x"b7",x"c8"),
    79 => (x"c1",x"87",x"c7",x"ff"),
    80 => (x"f0",x"c0",x"87",x"ce"),
    81 => (x"87",x"e6",x"c1",x"49"),
    82 => (x"c3",x"c1",x"84",x"c1"),
    83 => (x"73",x"83",x"c4",x"87"),
    84 => (x"6a",x"8a",x"c4",x"4a"),
    85 => (x"87",x"f1",x"c1",x"49"),
    86 => (x"4c",x"a4",x"49",x"70"),
    87 => (x"c4",x"87",x"f1",x"c0"),
    88 => (x"78",x"c1",x"48",x"a6"),
    89 => (x"c4",x"87",x"e9",x"c0"),
    90 => (x"c4",x"4a",x"73",x"83"),
    91 => (x"c0",x"49",x"6a",x"8a"),
    92 => (x"84",x"c1",x"87",x"fc"),
    93 => (x"49",x"6e",x"87",x"da"),
    94 => (x"d3",x"87",x"f3",x"c0"),
    95 => (x"c0",x"48",x"6e",x"87"),
    96 => (x"c7",x"05",x"a8",x"e5"),
    97 => (x"48",x"a6",x"c4",x"87"),
    98 => (x"87",x"c4",x"78",x"c1"),
    99 => (x"87",x"de",x"49",x"6e"),
   100 => (x"49",x"66",x"e0",x"c0"),
   101 => (x"c0",x"80",x"c1",x"48"),
   102 => (x"11",x"58",x"a6",x"e4"),
   103 => (x"fc",x"05",x"6e",x"7e"),
   104 => (x"48",x"74",x"87",x"cf"),
   105 => (x"4d",x"26",x"8e",x"f0"),
   106 => (x"4b",x"26",x"4c",x"26"),
   107 => (x"fc",x"1e",x"4f",x"26"),
   108 => (x"ff",x"4a",x"71",x"86"),
   109 => (x"48",x"69",x"49",x"c0"),
   110 => (x"70",x"98",x"c0",x"c4"),
   111 => (x"02",x"98",x"48",x"7e"),
   112 => (x"79",x"72",x"87",x"f4"),
   113 => (x"26",x"8e",x"fc",x"48"),
   114 => (x"5b",x"5e",x"0e",x"4f"),
   115 => (x"4b",x"71",x"0e",x"5c"),
   116 => (x"4a",x"13",x"4c",x"c0"),
   117 => (x"87",x"cd",x"02",x"9a"),
   118 => (x"d1",x"ff",x"49",x"72"),
   119 => (x"13",x"84",x"c1",x"87"),
   120 => (x"f3",x"05",x"9a",x"4a"),
   121 => (x"26",x"48",x"74",x"87"),
   122 => (x"26",x"4b",x"26",x"4c"),
   123 => (x"1e",x"72",x"1e",x"4f"),
   124 => (x"48",x"12",x"1e",x"73"),
   125 => (x"87",x"ca",x"02",x"11"),
   126 => (x"98",x"df",x"c3",x"4b"),
   127 => (x"02",x"88",x"73",x"9b"),
   128 => (x"4b",x"26",x"87",x"f0"),
   129 => (x"4f",x"26",x"4a",x"26"),
   130 => (x"72",x"1e",x"73",x"1e"),
   131 => (x"04",x"8b",x"c1",x"1e"),
   132 => (x"48",x"12",x"87",x"ca"),
   133 => (x"87",x"c4",x"02",x"11"),
   134 => (x"87",x"f1",x"02",x"88"),
   135 => (x"4b",x"26",x"4a",x"26"),
   136 => (x"73",x"1e",x"4f",x"26"),
   137 => (x"a9",x"73",x"81",x"48"),
   138 => (x"12",x"87",x"c5",x"02"),
   139 => (x"87",x"f6",x"05",x"53"),
   140 => (x"73",x"1e",x"4f",x"26"),
   141 => (x"c8",x"4a",x"71",x"1e"),
   142 => (x"c1",x"49",x"4b",x"66"),
   143 => (x"02",x"99",x"71",x"8b"),
   144 => (x"48",x"12",x"87",x"cf"),
   145 => (x"78",x"08",x"d4",x"ff"),
   146 => (x"8b",x"c1",x"49",x"73"),
   147 => (x"f1",x"05",x"99",x"71"),
   148 => (x"26",x"4b",x"26",x"87"),
   149 => (x"5b",x"5e",x"0e",x"4f"),
   150 => (x"4a",x"71",x"0e",x"5c"),
   151 => (x"cc",x"4c",x"d4",x"ff"),
   152 => (x"c1",x"49",x"4b",x"66"),
   153 => (x"02",x"99",x"71",x"8b"),
   154 => (x"ff",x"c3",x"87",x"ce"),
   155 => (x"73",x"52",x"6c",x"7c"),
   156 => (x"71",x"8b",x"c1",x"49"),
   157 => (x"87",x"f2",x"05",x"99"),
   158 => (x"4b",x"26",x"4c",x"26"),
   159 => (x"73",x"1e",x"4f",x"26"),
   160 => (x"4b",x"d4",x"ff",x"1e"),
   161 => (x"6b",x"7b",x"ff",x"c3"),
   162 => (x"7b",x"ff",x"c3",x"4a"),
   163 => (x"32",x"c8",x"49",x"6b"),
   164 => (x"ff",x"c3",x"b1",x"72"),
   165 => (x"c8",x"4a",x"6b",x"7b"),
   166 => (x"c3",x"b2",x"71",x"31"),
   167 => (x"49",x"6b",x"7b",x"ff"),
   168 => (x"b1",x"72",x"32",x"c8"),
   169 => (x"4b",x"26",x"48",x"71"),
   170 => (x"5e",x"0e",x"4f",x"26"),
   171 => (x"0e",x"5d",x"5c",x"5b"),
   172 => (x"d4",x"ff",x"4d",x"71"),
   173 => (x"c3",x"48",x"75",x"4c"),
   174 => (x"7c",x"70",x"98",x"ff"),
   175 => (x"bf",x"cc",x"e6",x"c2"),
   176 => (x"d0",x"87",x"c8",x"05"),
   177 => (x"30",x"c9",x"48",x"66"),
   178 => (x"d0",x"58",x"a6",x"d4"),
   179 => (x"29",x"d8",x"49",x"66"),
   180 => (x"ff",x"c3",x"48",x"71"),
   181 => (x"d0",x"7c",x"70",x"98"),
   182 => (x"29",x"d0",x"49",x"66"),
   183 => (x"ff",x"c3",x"48",x"71"),
   184 => (x"d0",x"7c",x"70",x"98"),
   185 => (x"29",x"c8",x"49",x"66"),
   186 => (x"ff",x"c3",x"48",x"71"),
   187 => (x"d0",x"7c",x"70",x"98"),
   188 => (x"ff",x"c3",x"48",x"66"),
   189 => (x"75",x"7c",x"70",x"98"),
   190 => (x"71",x"29",x"d0",x"49"),
   191 => (x"98",x"ff",x"c3",x"48"),
   192 => (x"4b",x"6c",x"7c",x"70"),
   193 => (x"4a",x"ff",x"f0",x"c9"),
   194 => (x"05",x"ab",x"ff",x"c3"),
   195 => (x"71",x"49",x"87",x"cf"),
   196 => (x"c1",x"4b",x"6c",x"7c"),
   197 => (x"87",x"c5",x"02",x"8a"),
   198 => (x"f2",x"02",x"ab",x"71"),
   199 => (x"26",x"48",x"73",x"87"),
   200 => (x"26",x"4c",x"26",x"4d"),
   201 => (x"1e",x"4f",x"26",x"4b"),
   202 => (x"d4",x"ff",x"49",x"c0"),
   203 => (x"78",x"ff",x"c3",x"48"),
   204 => (x"c8",x"c3",x"81",x"c1"),
   205 => (x"f1",x"04",x"a9",x"b7"),
   206 => (x"0e",x"4f",x"26",x"87"),
   207 => (x"5d",x"5c",x"5b",x"5e"),
   208 => (x"f0",x"ff",x"c0",x"0e"),
   209 => (x"c1",x"4d",x"f7",x"c1"),
   210 => (x"c0",x"c0",x"c0",x"c0"),
   211 => (x"d6",x"ff",x"4b",x"c0"),
   212 => (x"df",x"f8",x"c4",x"87"),
   213 => (x"75",x"1e",x"c0",x"4c"),
   214 => (x"87",x"ce",x"fd",x"49"),
   215 => (x"a8",x"c1",x"86",x"c4"),
   216 => (x"87",x"e5",x"c0",x"05"),
   217 => (x"c3",x"48",x"d4",x"ff"),
   218 => (x"1e",x"73",x"78",x"ff"),
   219 => (x"c1",x"f0",x"e1",x"c0"),
   220 => (x"f5",x"fc",x"49",x"e9"),
   221 => (x"70",x"86",x"c4",x"87"),
   222 => (x"87",x"ca",x"05",x"98"),
   223 => (x"c3",x"48",x"d4",x"ff"),
   224 => (x"48",x"c1",x"78",x"ff"),
   225 => (x"de",x"fe",x"87",x"cb"),
   226 => (x"05",x"8c",x"c1",x"87"),
   227 => (x"c0",x"87",x"c6",x"ff"),
   228 => (x"26",x"4d",x"26",x"48"),
   229 => (x"26",x"4b",x"26",x"4c"),
   230 => (x"5b",x"5e",x"0e",x"4f"),
   231 => (x"ff",x"c0",x"0e",x"5c"),
   232 => (x"4c",x"c1",x"c1",x"f0"),
   233 => (x"c3",x"48",x"d4",x"ff"),
   234 => (x"dc",x"cf",x"78",x"ff"),
   235 => (x"87",x"d9",x"f8",x"49"),
   236 => (x"1e",x"c0",x"4b",x"d3"),
   237 => (x"f1",x"fb",x"49",x"74"),
   238 => (x"70",x"86",x"c4",x"87"),
   239 => (x"87",x"ca",x"05",x"98"),
   240 => (x"c3",x"48",x"d4",x"ff"),
   241 => (x"48",x"c1",x"78",x"ff"),
   242 => (x"da",x"fd",x"87",x"cb"),
   243 => (x"05",x"8b",x"c1",x"87"),
   244 => (x"c0",x"87",x"df",x"ff"),
   245 => (x"26",x"4c",x"26",x"48"),
   246 => (x"00",x"4f",x"26",x"4b"),
   247 => (x"00",x"44",x"4d",x"43"),
   248 => (x"43",x"48",x"44",x"53"),
   249 => (x"69",x"61",x"66",x"20"),
   250 => (x"00",x"0a",x"21",x"6c"),
   251 => (x"52",x"52",x"45",x"49"),
   252 => (x"00",x"00",x"00",x"00"),
   253 => (x"00",x"49",x"50",x"53"),
   254 => (x"74",x"69",x"72",x"57"),
   255 => (x"61",x"66",x"20",x"65"),
   256 => (x"64",x"65",x"6c",x"69"),
   257 => (x"5e",x"0e",x"00",x"0a"),
   258 => (x"0e",x"5d",x"5c",x"5b"),
   259 => (x"ff",x"4d",x"ff",x"c3"),
   260 => (x"d2",x"fc",x"4b",x"d4"),
   261 => (x"1e",x"ea",x"c6",x"87"),
   262 => (x"c1",x"f0",x"e1",x"c0"),
   263 => (x"c9",x"fa",x"49",x"c8"),
   264 => (x"c1",x"86",x"c4",x"87"),
   265 => (x"87",x"c8",x"02",x"a8"),
   266 => (x"c0",x"87",x"ee",x"fd"),
   267 => (x"87",x"e8",x"c1",x"48"),
   268 => (x"70",x"87",x"cb",x"f9"),
   269 => (x"ff",x"ff",x"cf",x"49"),
   270 => (x"a9",x"ea",x"c6",x"99"),
   271 => (x"fd",x"87",x"c8",x"02"),
   272 => (x"48",x"c0",x"87",x"d7"),
   273 => (x"75",x"87",x"d1",x"c1"),
   274 => (x"4c",x"f1",x"c0",x"7b"),
   275 => (x"70",x"87",x"ec",x"fb"),
   276 => (x"ec",x"c0",x"02",x"98"),
   277 => (x"c0",x"1e",x"c0",x"87"),
   278 => (x"fa",x"c1",x"f0",x"ff"),
   279 => (x"87",x"ca",x"f9",x"49"),
   280 => (x"98",x"70",x"86",x"c4"),
   281 => (x"75",x"87",x"da",x"05"),
   282 => (x"75",x"49",x"6b",x"7b"),
   283 => (x"75",x"7b",x"75",x"7b"),
   284 => (x"c1",x"7b",x"75",x"7b"),
   285 => (x"c4",x"02",x"99",x"c0"),
   286 => (x"db",x"48",x"c1",x"87"),
   287 => (x"d7",x"48",x"c0",x"87"),
   288 => (x"05",x"ac",x"c2",x"87"),
   289 => (x"e0",x"cf",x"87",x"ca"),
   290 => (x"87",x"fd",x"f4",x"49"),
   291 => (x"87",x"c8",x"48",x"c0"),
   292 => (x"fe",x"05",x"8c",x"c1"),
   293 => (x"48",x"c0",x"87",x"f6"),
   294 => (x"4c",x"26",x"4d",x"26"),
   295 => (x"4f",x"26",x"4b",x"26"),
   296 => (x"5c",x"5b",x"5e",x"0e"),
   297 => (x"d0",x"ff",x"0e",x"5d"),
   298 => (x"d0",x"e5",x"c0",x"4d"),
   299 => (x"c2",x"4c",x"c0",x"c1"),
   300 => (x"c1",x"48",x"cc",x"e6"),
   301 => (x"49",x"f4",x"cf",x"78"),
   302 => (x"c7",x"87",x"ce",x"f4"),
   303 => (x"f9",x"7d",x"c2",x"4b"),
   304 => (x"7d",x"c3",x"87",x"e5"),
   305 => (x"49",x"74",x"1e",x"c0"),
   306 => (x"c4",x"87",x"df",x"f7"),
   307 => (x"05",x"a8",x"c1",x"86"),
   308 => (x"c2",x"4b",x"87",x"c1"),
   309 => (x"87",x"cb",x"05",x"ab"),
   310 => (x"f3",x"49",x"ec",x"cf"),
   311 => (x"48",x"c0",x"87",x"eb"),
   312 => (x"c1",x"87",x"f6",x"c0"),
   313 => (x"d4",x"ff",x"05",x"8b"),
   314 => (x"87",x"da",x"fc",x"87"),
   315 => (x"58",x"d0",x"e6",x"c2"),
   316 => (x"cd",x"05",x"98",x"70"),
   317 => (x"c0",x"1e",x"c1",x"87"),
   318 => (x"d0",x"c1",x"f0",x"ff"),
   319 => (x"87",x"ea",x"f6",x"49"),
   320 => (x"d4",x"ff",x"86",x"c4"),
   321 => (x"78",x"ff",x"c3",x"48"),
   322 => (x"c2",x"87",x"ee",x"c4"),
   323 => (x"c2",x"58",x"d4",x"e6"),
   324 => (x"48",x"d4",x"ff",x"7d"),
   325 => (x"c1",x"78",x"ff",x"c3"),
   326 => (x"26",x"4d",x"26",x"48"),
   327 => (x"26",x"4b",x"26",x"4c"),
   328 => (x"5b",x"5e",x"0e",x"4f"),
   329 => (x"71",x"0e",x"5d",x"5c"),
   330 => (x"4c",x"ff",x"c3",x"4d"),
   331 => (x"74",x"4b",x"d4",x"ff"),
   332 => (x"48",x"d0",x"ff",x"7b"),
   333 => (x"74",x"78",x"c3",x"c4"),
   334 => (x"c0",x"1e",x"75",x"7b"),
   335 => (x"d8",x"c1",x"f0",x"ff"),
   336 => (x"87",x"e6",x"f5",x"49"),
   337 => (x"98",x"70",x"86",x"c4"),
   338 => (x"cf",x"87",x"cb",x"02"),
   339 => (x"f8",x"f1",x"49",x"f8"),
   340 => (x"c0",x"48",x"c1",x"87"),
   341 => (x"7b",x"74",x"87",x"ee"),
   342 => (x"c8",x"7b",x"fe",x"c3"),
   343 => (x"66",x"d4",x"1e",x"c0"),
   344 => (x"87",x"ce",x"f3",x"49"),
   345 => (x"7b",x"74",x"86",x"c4"),
   346 => (x"7b",x"74",x"7b",x"74"),
   347 => (x"4a",x"e0",x"da",x"d8"),
   348 => (x"05",x"6b",x"7b",x"74"),
   349 => (x"8a",x"c1",x"87",x"c5"),
   350 => (x"74",x"87",x"f5",x"05"),
   351 => (x"48",x"d0",x"ff",x"7b"),
   352 => (x"48",x"c0",x"78",x"c2"),
   353 => (x"4c",x"26",x"4d",x"26"),
   354 => (x"4f",x"26",x"4b",x"26"),
   355 => (x"5c",x"5b",x"5e",x"0e"),
   356 => (x"86",x"fc",x"0e",x"5d"),
   357 => (x"d4",x"ff",x"4b",x"71"),
   358 => (x"c5",x"7e",x"c0",x"4c"),
   359 => (x"4a",x"df",x"cd",x"ee"),
   360 => (x"6c",x"7c",x"ff",x"c3"),
   361 => (x"a8",x"fe",x"c3",x"48"),
   362 => (x"87",x"f8",x"c0",x"05"),
   363 => (x"9b",x"73",x"4d",x"74"),
   364 => (x"d4",x"87",x"cc",x"02"),
   365 => (x"49",x"73",x"1e",x"66"),
   366 => (x"c4",x"87",x"da",x"f2"),
   367 => (x"ff",x"87",x"d4",x"86"),
   368 => (x"d1",x"c4",x"48",x"d0"),
   369 => (x"4a",x"66",x"d4",x"78"),
   370 => (x"c1",x"7d",x"ff",x"c3"),
   371 => (x"87",x"f8",x"05",x"8a"),
   372 => (x"c3",x"5a",x"a6",x"d8"),
   373 => (x"73",x"7c",x"7c",x"ff"),
   374 => (x"87",x"c5",x"05",x"9b"),
   375 => (x"d0",x"48",x"d0",x"ff"),
   376 => (x"7e",x"4a",x"c1",x"78"),
   377 => (x"fe",x"05",x"8a",x"c1"),
   378 => (x"48",x"6e",x"87",x"f6"),
   379 => (x"4d",x"26",x"8e",x"fc"),
   380 => (x"4b",x"26",x"4c",x"26"),
   381 => (x"73",x"1e",x"4f",x"26"),
   382 => (x"c0",x"4a",x"71",x"1e"),
   383 => (x"48",x"d4",x"ff",x"4b"),
   384 => (x"ff",x"78",x"ff",x"c3"),
   385 => (x"c3",x"c4",x"48",x"d0"),
   386 => (x"48",x"d4",x"ff",x"78"),
   387 => (x"72",x"78",x"ff",x"c3"),
   388 => (x"f0",x"ff",x"c0",x"1e"),
   389 => (x"f2",x"49",x"d1",x"c1"),
   390 => (x"86",x"c4",x"87",x"d0"),
   391 => (x"d2",x"05",x"98",x"70"),
   392 => (x"1e",x"c0",x"c8",x"87"),
   393 => (x"fd",x"49",x"66",x"cc"),
   394 => (x"86",x"c4",x"87",x"e2"),
   395 => (x"d0",x"ff",x"4b",x"70"),
   396 => (x"73",x"78",x"c2",x"48"),
   397 => (x"26",x"4b",x"26",x"48"),
   398 => (x"5b",x"5e",x"0e",x"4f"),
   399 => (x"c0",x"0e",x"5d",x"5c"),
   400 => (x"f0",x"ff",x"c0",x"1e"),
   401 => (x"f1",x"49",x"c9",x"c1"),
   402 => (x"1e",x"d2",x"87",x"e0"),
   403 => (x"49",x"dc",x"e6",x"c2"),
   404 => (x"c8",x"87",x"f9",x"fc"),
   405 => (x"c1",x"4c",x"c0",x"86"),
   406 => (x"ac",x"b7",x"d2",x"84"),
   407 => (x"c2",x"87",x"f8",x"04"),
   408 => (x"bf",x"97",x"dc",x"e6"),
   409 => (x"99",x"c0",x"c3",x"49"),
   410 => (x"05",x"a9",x"c0",x"c1"),
   411 => (x"c2",x"87",x"e7",x"c0"),
   412 => (x"bf",x"97",x"e3",x"e6"),
   413 => (x"c2",x"31",x"d0",x"49"),
   414 => (x"bf",x"97",x"e4",x"e6"),
   415 => (x"72",x"32",x"c8",x"4a"),
   416 => (x"e5",x"e6",x"c2",x"b1"),
   417 => (x"b1",x"4a",x"bf",x"97"),
   418 => (x"ff",x"cf",x"4c",x"71"),
   419 => (x"c1",x"9c",x"ff",x"ff"),
   420 => (x"c1",x"34",x"ca",x"84"),
   421 => (x"e6",x"c2",x"87",x"e7"),
   422 => (x"49",x"bf",x"97",x"e5"),
   423 => (x"99",x"c6",x"31",x"c1"),
   424 => (x"97",x"e6",x"e6",x"c2"),
   425 => (x"b7",x"c7",x"4a",x"bf"),
   426 => (x"c2",x"b1",x"72",x"2a"),
   427 => (x"bf",x"97",x"e1",x"e6"),
   428 => (x"9d",x"cf",x"4d",x"4a"),
   429 => (x"97",x"e2",x"e6",x"c2"),
   430 => (x"9a",x"c3",x"4a",x"bf"),
   431 => (x"e6",x"c2",x"32",x"ca"),
   432 => (x"4b",x"bf",x"97",x"e3"),
   433 => (x"b2",x"73",x"33",x"c2"),
   434 => (x"97",x"e4",x"e6",x"c2"),
   435 => (x"c0",x"c3",x"4b",x"bf"),
   436 => (x"2b",x"b7",x"c6",x"9b"),
   437 => (x"81",x"c2",x"b2",x"73"),
   438 => (x"30",x"71",x"48",x"c1"),
   439 => (x"48",x"c1",x"49",x"70"),
   440 => (x"4d",x"70",x"30",x"75"),
   441 => (x"84",x"c1",x"4c",x"72"),
   442 => (x"c0",x"c8",x"94",x"71"),
   443 => (x"cc",x"06",x"ad",x"b7"),
   444 => (x"b7",x"34",x"c1",x"87"),
   445 => (x"b7",x"c0",x"c8",x"2d"),
   446 => (x"f4",x"ff",x"01",x"ad"),
   447 => (x"26",x"48",x"74",x"87"),
   448 => (x"26",x"4c",x"26",x"4d"),
   449 => (x"0e",x"4f",x"26",x"4b"),
   450 => (x"5d",x"5c",x"5b",x"5e"),
   451 => (x"c2",x"86",x"fc",x"0e"),
   452 => (x"c0",x"48",x"c4",x"ef"),
   453 => (x"fc",x"e6",x"c2",x"78"),
   454 => (x"fb",x"49",x"c0",x"1e"),
   455 => (x"86",x"c4",x"87",x"d8"),
   456 => (x"c5",x"05",x"98",x"70"),
   457 => (x"c9",x"48",x"c0",x"87"),
   458 => (x"4d",x"c0",x"87",x"d5"),
   459 => (x"48",x"c0",x"f4",x"c2"),
   460 => (x"e7",x"c2",x"78",x"c1"),
   461 => (x"e6",x"c0",x"4a",x"f2"),
   462 => (x"4b",x"c8",x"49",x"d8"),
   463 => (x"70",x"87",x"c9",x"eb"),
   464 => (x"87",x"c6",x"05",x"98"),
   465 => (x"48",x"c0",x"f4",x"c2"),
   466 => (x"e8",x"c2",x"78",x"c0"),
   467 => (x"e6",x"c0",x"4a",x"ce"),
   468 => (x"4b",x"c8",x"49",x"e4"),
   469 => (x"70",x"87",x"f1",x"ea"),
   470 => (x"87",x"c6",x"05",x"98"),
   471 => (x"48",x"c0",x"f4",x"c2"),
   472 => (x"f4",x"c2",x"78",x"c0"),
   473 => (x"c0",x"02",x"bf",x"c0"),
   474 => (x"ee",x"c2",x"87",x"fe"),
   475 => (x"c2",x"4d",x"bf",x"c2"),
   476 => (x"bf",x"9f",x"fa",x"ee"),
   477 => (x"c5",x"48",x"6e",x"7e"),
   478 => (x"05",x"a8",x"ea",x"d6"),
   479 => (x"ee",x"c2",x"87",x"c7"),
   480 => (x"ce",x"4d",x"bf",x"c2"),
   481 => (x"ca",x"48",x"6e",x"87"),
   482 => (x"02",x"a8",x"d5",x"e9"),
   483 => (x"48",x"c0",x"87",x"c5"),
   484 => (x"c2",x"87",x"ec",x"c7"),
   485 => (x"75",x"1e",x"fc",x"e6"),
   486 => (x"87",x"da",x"f9",x"49"),
   487 => (x"98",x"70",x"86",x"c4"),
   488 => (x"c0",x"87",x"c5",x"05"),
   489 => (x"87",x"d7",x"c7",x"48"),
   490 => (x"4a",x"ce",x"e8",x"c2"),
   491 => (x"49",x"f0",x"e6",x"c0"),
   492 => (x"d3",x"e9",x"4b",x"c8"),
   493 => (x"05",x"98",x"70",x"87"),
   494 => (x"c2",x"87",x"c8",x"c0"),
   495 => (x"c1",x"48",x"c4",x"ef"),
   496 => (x"c2",x"87",x"d8",x"78"),
   497 => (x"c0",x"4a",x"f2",x"e7"),
   498 => (x"c8",x"49",x"fc",x"e6"),
   499 => (x"87",x"f8",x"e8",x"4b"),
   500 => (x"c0",x"02",x"98",x"70"),
   501 => (x"48",x"c0",x"87",x"c5"),
   502 => (x"c2",x"87",x"e4",x"c6"),
   503 => (x"bf",x"97",x"fa",x"ee"),
   504 => (x"a9",x"d5",x"c1",x"49"),
   505 => (x"87",x"cd",x"c0",x"05"),
   506 => (x"97",x"fb",x"ee",x"c2"),
   507 => (x"ea",x"c2",x"49",x"bf"),
   508 => (x"c5",x"c0",x"02",x"a9"),
   509 => (x"c6",x"48",x"c0",x"87"),
   510 => (x"e6",x"c2",x"87",x"c5"),
   511 => (x"7e",x"bf",x"97",x"fc"),
   512 => (x"e9",x"c3",x"48",x"6e"),
   513 => (x"ce",x"c0",x"02",x"a8"),
   514 => (x"c3",x"48",x"6e",x"87"),
   515 => (x"c0",x"02",x"a8",x"eb"),
   516 => (x"48",x"c0",x"87",x"c5"),
   517 => (x"c2",x"87",x"e8",x"c5"),
   518 => (x"bf",x"97",x"c7",x"e7"),
   519 => (x"c0",x"05",x"99",x"49"),
   520 => (x"e7",x"c2",x"87",x"cc"),
   521 => (x"49",x"bf",x"97",x"c8"),
   522 => (x"c0",x"02",x"a9",x"c2"),
   523 => (x"48",x"c0",x"87",x"c5"),
   524 => (x"c2",x"87",x"cc",x"c5"),
   525 => (x"bf",x"97",x"c9",x"e7"),
   526 => (x"c0",x"ef",x"c2",x"48"),
   527 => (x"48",x"4c",x"70",x"58"),
   528 => (x"ef",x"c2",x"88",x"c1"),
   529 => (x"e7",x"c2",x"58",x"c4"),
   530 => (x"49",x"bf",x"97",x"ca"),
   531 => (x"e7",x"c2",x"81",x"75"),
   532 => (x"4a",x"bf",x"97",x"cb"),
   533 => (x"a1",x"72",x"32",x"c8"),
   534 => (x"dc",x"f3",x"c2",x"7e"),
   535 => (x"c2",x"78",x"6e",x"48"),
   536 => (x"bf",x"97",x"cc",x"e7"),
   537 => (x"f4",x"f3",x"c2",x"48"),
   538 => (x"c4",x"ef",x"c2",x"58"),
   539 => (x"d3",x"c2",x"02",x"bf"),
   540 => (x"ce",x"e8",x"c2",x"87"),
   541 => (x"cc",x"e6",x"c0",x"4a"),
   542 => (x"e6",x"4b",x"c8",x"49"),
   543 => (x"98",x"70",x"87",x"ca"),
   544 => (x"87",x"c5",x"c0",x"02"),
   545 => (x"f6",x"c3",x"48",x"c0"),
   546 => (x"fc",x"ee",x"c2",x"87"),
   547 => (x"f3",x"c2",x"4c",x"bf"),
   548 => (x"e7",x"c2",x"5c",x"f0"),
   549 => (x"49",x"bf",x"97",x"e1"),
   550 => (x"e7",x"c2",x"31",x"c8"),
   551 => (x"4a",x"bf",x"97",x"e0"),
   552 => (x"e7",x"c2",x"49",x"a1"),
   553 => (x"4a",x"bf",x"97",x"e2"),
   554 => (x"a1",x"72",x"32",x"d0"),
   555 => (x"e3",x"e7",x"c2",x"49"),
   556 => (x"d8",x"4a",x"bf",x"97"),
   557 => (x"49",x"a1",x"72",x"32"),
   558 => (x"59",x"f8",x"f3",x"c2"),
   559 => (x"bf",x"f0",x"f3",x"c2"),
   560 => (x"dc",x"f3",x"c2",x"91"),
   561 => (x"f3",x"c2",x"81",x"bf"),
   562 => (x"e7",x"c2",x"59",x"e4"),
   563 => (x"4a",x"bf",x"97",x"e9"),
   564 => (x"e7",x"c2",x"32",x"c8"),
   565 => (x"4b",x"bf",x"97",x"e8"),
   566 => (x"e7",x"c2",x"4a",x"a2"),
   567 => (x"4b",x"bf",x"97",x"ea"),
   568 => (x"a2",x"73",x"33",x"d0"),
   569 => (x"eb",x"e7",x"c2",x"4a"),
   570 => (x"cf",x"4b",x"bf",x"97"),
   571 => (x"73",x"33",x"d8",x"9b"),
   572 => (x"f3",x"c2",x"4a",x"a2"),
   573 => (x"8a",x"c2",x"5a",x"e8"),
   574 => (x"f3",x"c2",x"92",x"74"),
   575 => (x"a1",x"72",x"48",x"e8"),
   576 => (x"87",x"c7",x"c1",x"78"),
   577 => (x"97",x"ce",x"e7",x"c2"),
   578 => (x"31",x"c8",x"49",x"bf"),
   579 => (x"97",x"cd",x"e7",x"c2"),
   580 => (x"49",x"a1",x"4a",x"bf"),
   581 => (x"ff",x"c7",x"31",x"c5"),
   582 => (x"c2",x"29",x"c9",x"81"),
   583 => (x"c2",x"59",x"f0",x"f3"),
   584 => (x"bf",x"97",x"d3",x"e7"),
   585 => (x"c2",x"32",x"c8",x"4a"),
   586 => (x"bf",x"97",x"d2",x"e7"),
   587 => (x"c2",x"4a",x"a2",x"4b"),
   588 => (x"c2",x"5a",x"f8",x"f3"),
   589 => (x"92",x"bf",x"f0",x"f3"),
   590 => (x"f3",x"c2",x"82",x"6e"),
   591 => (x"f3",x"c2",x"5a",x"ec"),
   592 => (x"78",x"c0",x"48",x"e4"),
   593 => (x"48",x"e0",x"f3",x"c2"),
   594 => (x"c2",x"78",x"a1",x"72"),
   595 => (x"c2",x"48",x"f8",x"f3"),
   596 => (x"78",x"bf",x"e4",x"f3"),
   597 => (x"48",x"fc",x"f3",x"c2"),
   598 => (x"bf",x"e8",x"f3",x"c2"),
   599 => (x"c4",x"ef",x"c2",x"78"),
   600 => (x"c9",x"c0",x"02",x"bf"),
   601 => (x"c4",x"48",x"74",x"87"),
   602 => (x"c0",x"7e",x"70",x"30"),
   603 => (x"f3",x"c2",x"87",x"c9"),
   604 => (x"c4",x"48",x"bf",x"ec"),
   605 => (x"c2",x"7e",x"70",x"30"),
   606 => (x"6e",x"48",x"c8",x"ef"),
   607 => (x"fc",x"48",x"c1",x"78"),
   608 => (x"26",x"4d",x"26",x"8e"),
   609 => (x"26",x"4b",x"26",x"4c"),
   610 => (x"00",x"00",x"00",x"4f"),
   611 => (x"33",x"54",x"41",x"46"),
   612 => (x"20",x"20",x"20",x"32"),
   613 => (x"00",x"00",x"00",x"00"),
   614 => (x"31",x"54",x"41",x"46"),
   615 => (x"20",x"20",x"20",x"36"),
   616 => (x"00",x"00",x"00",x"00"),
   617 => (x"33",x"54",x"41",x"46"),
   618 => (x"20",x"20",x"20",x"32"),
   619 => (x"00",x"00",x"00",x"00"),
   620 => (x"33",x"54",x"41",x"46"),
   621 => (x"20",x"20",x"20",x"32"),
   622 => (x"00",x"00",x"00",x"00"),
   623 => (x"31",x"54",x"41",x"46"),
   624 => (x"20",x"20",x"20",x"36"),
   625 => (x"5b",x"5e",x"0e",x"00"),
   626 => (x"71",x"0e",x"5d",x"5c"),
   627 => (x"c4",x"ef",x"c2",x"4a"),
   628 => (x"87",x"cb",x"02",x"bf"),
   629 => (x"2b",x"c7",x"4b",x"72"),
   630 => (x"ff",x"c1",x"4d",x"72"),
   631 => (x"72",x"87",x"c9",x"9d"),
   632 => (x"72",x"2b",x"c8",x"4b"),
   633 => (x"9d",x"ff",x"c3",x"4d"),
   634 => (x"bf",x"dc",x"f3",x"c2"),
   635 => (x"d0",x"fe",x"c0",x"83"),
   636 => (x"d9",x"02",x"ab",x"bf"),
   637 => (x"d4",x"fe",x"c0",x"87"),
   638 => (x"fc",x"e6",x"c2",x"5b"),
   639 => (x"ef",x"49",x"73",x"1e"),
   640 => (x"86",x"c4",x"87",x"f4"),
   641 => (x"c5",x"05",x"98",x"70"),
   642 => (x"c0",x"48",x"c0",x"87"),
   643 => (x"ef",x"c2",x"87",x"e6"),
   644 => (x"d2",x"02",x"bf",x"c4"),
   645 => (x"c4",x"49",x"75",x"87"),
   646 => (x"fc",x"e6",x"c2",x"91"),
   647 => (x"cf",x"4c",x"69",x"81"),
   648 => (x"ff",x"ff",x"ff",x"ff"),
   649 => (x"75",x"87",x"cb",x"9c"),
   650 => (x"c2",x"91",x"c2",x"49"),
   651 => (x"9f",x"81",x"fc",x"e6"),
   652 => (x"48",x"74",x"4c",x"69"),
   653 => (x"4c",x"26",x"4d",x"26"),
   654 => (x"4f",x"26",x"4b",x"26"),
   655 => (x"5c",x"5b",x"5e",x"0e"),
   656 => (x"86",x"f4",x"0e",x"5d"),
   657 => (x"c4",x"59",x"a6",x"c8"),
   658 => (x"80",x"c8",x"48",x"66"),
   659 => (x"48",x"6e",x"7e",x"70"),
   660 => (x"c1",x"1e",x"78",x"c0"),
   661 => (x"87",x"fd",x"cc",x"49"),
   662 => (x"4c",x"70",x"86",x"c4"),
   663 => (x"fc",x"c0",x"02",x"9c"),
   664 => (x"cc",x"ef",x"c2",x"87"),
   665 => (x"49",x"66",x"dc",x"4a"),
   666 => (x"87",x"c1",x"de",x"ff"),
   667 => (x"c0",x"02",x"98",x"70"),
   668 => (x"4a",x"74",x"87",x"eb"),
   669 => (x"cb",x"49",x"66",x"dc"),
   670 => (x"cb",x"de",x"ff",x"4b"),
   671 => (x"02",x"98",x"70",x"87"),
   672 => (x"1e",x"c0",x"87",x"db"),
   673 => (x"c4",x"02",x"9c",x"74"),
   674 => (x"c2",x"4d",x"c0",x"87"),
   675 => (x"75",x"4d",x"c1",x"87"),
   676 => (x"87",x"c1",x"cc",x"49"),
   677 => (x"4c",x"70",x"86",x"c4"),
   678 => (x"c4",x"ff",x"05",x"9c"),
   679 => (x"02",x"9c",x"74",x"87"),
   680 => (x"dc",x"87",x"f4",x"c1"),
   681 => (x"48",x"6e",x"49",x"a4"),
   682 => (x"a4",x"da",x"78",x"69"),
   683 => (x"4d",x"66",x"c4",x"49"),
   684 => (x"69",x"9f",x"85",x"c4"),
   685 => (x"c4",x"ef",x"c2",x"7d"),
   686 => (x"87",x"d2",x"02",x"bf"),
   687 => (x"9f",x"49",x"a4",x"d4"),
   688 => (x"ff",x"c0",x"49",x"69"),
   689 => (x"48",x"71",x"99",x"ff"),
   690 => (x"7e",x"70",x"30",x"d0"),
   691 => (x"7e",x"c0",x"87",x"c2"),
   692 => (x"6d",x"48",x"49",x"6e"),
   693 => (x"c4",x"7d",x"70",x"80"),
   694 => (x"78",x"c0",x"48",x"66"),
   695 => (x"cc",x"49",x"66",x"c4"),
   696 => (x"c4",x"79",x"6d",x"81"),
   697 => (x"81",x"d0",x"49",x"66"),
   698 => (x"a6",x"c8",x"79",x"c0"),
   699 => (x"c8",x"78",x"c0",x"48"),
   700 => (x"66",x"c4",x"4c",x"66"),
   701 => (x"74",x"82",x"d4",x"4a"),
   702 => (x"72",x"91",x"c8",x"49"),
   703 => (x"41",x"c0",x"49",x"a1"),
   704 => (x"84",x"c1",x"79",x"6d"),
   705 => (x"04",x"ac",x"b7",x"c6"),
   706 => (x"c4",x"87",x"e7",x"ff"),
   707 => (x"c4",x"c1",x"49",x"66"),
   708 => (x"c1",x"79",x"c0",x"81"),
   709 => (x"c0",x"87",x"c2",x"48"),
   710 => (x"26",x"8e",x"f4",x"48"),
   711 => (x"26",x"4c",x"26",x"4d"),
   712 => (x"0e",x"4f",x"26",x"4b"),
   713 => (x"5d",x"5c",x"5b",x"5e"),
   714 => (x"d0",x"4c",x"71",x"0e"),
   715 => (x"49",x"6c",x"4d",x"66"),
   716 => (x"c2",x"b9",x"75",x"85"),
   717 => (x"4a",x"bf",x"c0",x"ef"),
   718 => (x"99",x"72",x"ba",x"ff"),
   719 => (x"c0",x"02",x"99",x"71"),
   720 => (x"a4",x"c4",x"87",x"e4"),
   721 => (x"f9",x"49",x"6b",x"4b"),
   722 => (x"7b",x"70",x"87",x"fb"),
   723 => (x"bf",x"fc",x"ee",x"c2"),
   724 => (x"71",x"81",x"6c",x"49"),
   725 => (x"c2",x"b9",x"75",x"7c"),
   726 => (x"4a",x"bf",x"c0",x"ef"),
   727 => (x"99",x"72",x"ba",x"ff"),
   728 => (x"ff",x"05",x"99",x"71"),
   729 => (x"7c",x"75",x"87",x"dc"),
   730 => (x"4c",x"26",x"4d",x"26"),
   731 => (x"4f",x"26",x"4b",x"26"),
   732 => (x"71",x"1e",x"73",x"1e"),
   733 => (x"e0",x"f3",x"c2",x"4b"),
   734 => (x"a3",x"c4",x"49",x"bf"),
   735 => (x"c2",x"4a",x"6a",x"4a"),
   736 => (x"fc",x"ee",x"c2",x"8a"),
   737 => (x"a1",x"72",x"92",x"bf"),
   738 => (x"c0",x"ef",x"c2",x"49"),
   739 => (x"9a",x"6b",x"4a",x"bf"),
   740 => (x"c0",x"49",x"a1",x"72"),
   741 => (x"c8",x"59",x"d4",x"fe"),
   742 => (x"e9",x"71",x"1e",x"66"),
   743 => (x"86",x"c4",x"87",x"d8"),
   744 => (x"c4",x"05",x"98",x"70"),
   745 => (x"c2",x"48",x"c0",x"87"),
   746 => (x"26",x"48",x"c1",x"87"),
   747 => (x"1e",x"4f",x"26",x"4b"),
   748 => (x"4b",x"71",x"1e",x"73"),
   749 => (x"bf",x"e0",x"f3",x"c2"),
   750 => (x"4a",x"a3",x"c4",x"49"),
   751 => (x"8a",x"c2",x"4a",x"6a"),
   752 => (x"bf",x"fc",x"ee",x"c2"),
   753 => (x"49",x"a1",x"72",x"92"),
   754 => (x"bf",x"c0",x"ef",x"c2"),
   755 => (x"72",x"9a",x"6b",x"4a"),
   756 => (x"fe",x"c0",x"49",x"a1"),
   757 => (x"66",x"c8",x"59",x"d4"),
   758 => (x"c4",x"e5",x"71",x"1e"),
   759 => (x"70",x"86",x"c4",x"87"),
   760 => (x"87",x"c4",x"05",x"98"),
   761 => (x"87",x"c2",x"48",x"c0"),
   762 => (x"4b",x"26",x"48",x"c1"),
   763 => (x"5e",x"0e",x"4f",x"26"),
   764 => (x"0e",x"5d",x"5c",x"5b"),
   765 => (x"4b",x"71",x"86",x"e4"),
   766 => (x"48",x"66",x"ec",x"c0"),
   767 => (x"a6",x"cc",x"28",x"c9"),
   768 => (x"c0",x"ef",x"c2",x"58"),
   769 => (x"b9",x"ff",x"49",x"bf"),
   770 => (x"66",x"c8",x"48",x"71"),
   771 => (x"58",x"a6",x"d4",x"98"),
   772 => (x"98",x"6b",x"48",x"71"),
   773 => (x"c4",x"58",x"a6",x"d0"),
   774 => (x"a6",x"c4",x"7e",x"a3"),
   775 => (x"78",x"bf",x"6e",x"48"),
   776 => (x"cc",x"48",x"66",x"d0"),
   777 => (x"c6",x"05",x"a8",x"66"),
   778 => (x"7b",x"66",x"c8",x"87"),
   779 => (x"d4",x"87",x"c6",x"c3"),
   780 => (x"ff",x"c1",x"48",x"a6"),
   781 => (x"ff",x"ff",x"ff",x"ff"),
   782 => (x"ff",x"80",x"c4",x"78"),
   783 => (x"d4",x"4a",x"c0",x"78"),
   784 => (x"49",x"72",x"4d",x"a3"),
   785 => (x"a1",x"75",x"91",x"c8"),
   786 => (x"4c",x"66",x"d0",x"49"),
   787 => (x"b7",x"c0",x"8c",x"69"),
   788 => (x"87",x"cd",x"04",x"ac"),
   789 => (x"ac",x"b7",x"66",x"d4"),
   790 => (x"dc",x"87",x"c6",x"03"),
   791 => (x"a6",x"d8",x"5a",x"a6"),
   792 => (x"c6",x"82",x"c1",x"5c"),
   793 => (x"ff",x"04",x"aa",x"b7"),
   794 => (x"66",x"d8",x"87",x"d5"),
   795 => (x"a8",x"b7",x"c0",x"48"),
   796 => (x"d8",x"87",x"d0",x"04"),
   797 => (x"91",x"c8",x"49",x"66"),
   798 => (x"21",x"49",x"a1",x"75"),
   799 => (x"69",x"48",x"6e",x"7b"),
   800 => (x"c0",x"87",x"c9",x"78"),
   801 => (x"49",x"a3",x"cc",x"7b"),
   802 => (x"78",x"69",x"48",x"6e"),
   803 => (x"6b",x"48",x"66",x"c8"),
   804 => (x"58",x"a6",x"cc",x"88"),
   805 => (x"bf",x"fc",x"ee",x"c2"),
   806 => (x"70",x"90",x"c8",x"48"),
   807 => (x"48",x"66",x"c8",x"7e"),
   808 => (x"c9",x"01",x"a8",x"6e"),
   809 => (x"48",x"66",x"c8",x"87"),
   810 => (x"c0",x"03",x"a8",x"6e"),
   811 => (x"c4",x"c1",x"87",x"fd"),
   812 => (x"bf",x"6e",x"7e",x"a3"),
   813 => (x"75",x"91",x"c8",x"49"),
   814 => (x"66",x"cc",x"49",x"a1"),
   815 => (x"49",x"bf",x"6e",x"79"),
   816 => (x"a1",x"75",x"91",x"c8"),
   817 => (x"66",x"81",x"c4",x"49"),
   818 => (x"48",x"a6",x"d0",x"79"),
   819 => (x"d0",x"78",x"bf",x"6e"),
   820 => (x"a8",x"c5",x"48",x"66"),
   821 => (x"c4",x"87",x"c7",x"05"),
   822 => (x"78",x"c0",x"48",x"a6"),
   823 => (x"66",x"d0",x"87",x"c8"),
   824 => (x"c8",x"80",x"c1",x"48"),
   825 => (x"48",x"6e",x"58",x"a6"),
   826 => (x"c8",x"78",x"66",x"c4"),
   827 => (x"49",x"73",x"1e",x"66"),
   828 => (x"c4",x"87",x"f0",x"f8"),
   829 => (x"fc",x"e6",x"c2",x"86"),
   830 => (x"f9",x"49",x"73",x"1e"),
   831 => (x"a3",x"d0",x"87",x"f2"),
   832 => (x"66",x"f0",x"c0",x"49"),
   833 => (x"26",x"8e",x"e0",x"79"),
   834 => (x"26",x"4c",x"26",x"4d"),
   835 => (x"0e",x"4f",x"26",x"4b"),
   836 => (x"0e",x"5c",x"5b",x"5e"),
   837 => (x"4b",x"c0",x"4a",x"71"),
   838 => (x"c0",x"02",x"9a",x"72"),
   839 => (x"a2",x"da",x"87",x"e0"),
   840 => (x"4b",x"69",x"9f",x"49"),
   841 => (x"bf",x"c4",x"ef",x"c2"),
   842 => (x"d4",x"87",x"cf",x"02"),
   843 => (x"69",x"9f",x"49",x"a2"),
   844 => (x"ff",x"c0",x"4c",x"49"),
   845 => (x"34",x"d0",x"9c",x"ff"),
   846 => (x"4c",x"c0",x"87",x"c2"),
   847 => (x"9b",x"73",x"b3",x"74"),
   848 => (x"4a",x"87",x"df",x"02"),
   849 => (x"ee",x"c2",x"8a",x"c2"),
   850 => (x"92",x"49",x"bf",x"fc"),
   851 => (x"bf",x"e0",x"f3",x"c2"),
   852 => (x"c2",x"80",x"72",x"48"),
   853 => (x"71",x"58",x"c0",x"f4"),
   854 => (x"c2",x"30",x"c4",x"48"),
   855 => (x"c0",x"58",x"cc",x"ef"),
   856 => (x"f3",x"c2",x"87",x"e9"),
   857 => (x"c2",x"4b",x"bf",x"e4"),
   858 => (x"c2",x"48",x"fc",x"f3"),
   859 => (x"78",x"bf",x"e8",x"f3"),
   860 => (x"bf",x"c4",x"ef",x"c2"),
   861 => (x"c2",x"87",x"c9",x"02"),
   862 => (x"49",x"bf",x"fc",x"ee"),
   863 => (x"87",x"c7",x"31",x"c4"),
   864 => (x"bf",x"ec",x"f3",x"c2"),
   865 => (x"c2",x"31",x"c4",x"49"),
   866 => (x"c2",x"59",x"cc",x"ef"),
   867 => (x"26",x"5b",x"fc",x"f3"),
   868 => (x"26",x"4b",x"26",x"4c"),
   869 => (x"5b",x"5e",x"0e",x"4f"),
   870 => (x"f0",x"0e",x"5d",x"5c"),
   871 => (x"59",x"a6",x"c8",x"86"),
   872 => (x"ff",x"ff",x"ff",x"cf"),
   873 => (x"7e",x"c0",x"4c",x"f8"),
   874 => (x"d8",x"02",x"66",x"c4"),
   875 => (x"f8",x"e6",x"c2",x"87"),
   876 => (x"c2",x"78",x"c0",x"48"),
   877 => (x"c2",x"48",x"f0",x"e6"),
   878 => (x"78",x"bf",x"fc",x"f3"),
   879 => (x"48",x"f4",x"e6",x"c2"),
   880 => (x"bf",x"f8",x"f3",x"c2"),
   881 => (x"d9",x"ef",x"c2",x"78"),
   882 => (x"c2",x"50",x"c0",x"48"),
   883 => (x"49",x"bf",x"c8",x"ef"),
   884 => (x"bf",x"f8",x"e6",x"c2"),
   885 => (x"03",x"aa",x"71",x"4a"),
   886 => (x"72",x"87",x"cc",x"c4"),
   887 => (x"05",x"99",x"cf",x"49"),
   888 => (x"c0",x"87",x"ea",x"c0"),
   889 => (x"c2",x"48",x"d0",x"fe"),
   890 => (x"78",x"bf",x"f0",x"e6"),
   891 => (x"1e",x"fc",x"e6",x"c2"),
   892 => (x"bf",x"f0",x"e6",x"c2"),
   893 => (x"f0",x"e6",x"c2",x"49"),
   894 => (x"78",x"a1",x"c1",x"48"),
   895 => (x"f5",x"df",x"ff",x"71"),
   896 => (x"c0",x"86",x"c4",x"87"),
   897 => (x"c2",x"48",x"cc",x"fe"),
   898 => (x"cc",x"78",x"fc",x"e6"),
   899 => (x"cc",x"fe",x"c0",x"87"),
   900 => (x"e0",x"c0",x"48",x"bf"),
   901 => (x"d0",x"fe",x"c0",x"80"),
   902 => (x"f8",x"e6",x"c2",x"58"),
   903 => (x"80",x"c1",x"48",x"bf"),
   904 => (x"58",x"fc",x"e6",x"c2"),
   905 => (x"00",x"0f",x"8c",x"27"),
   906 => (x"bf",x"97",x"bf",x"00"),
   907 => (x"c2",x"02",x"9d",x"4d"),
   908 => (x"e5",x"c3",x"87",x"e5"),
   909 => (x"de",x"c2",x"02",x"ad"),
   910 => (x"cc",x"fe",x"c0",x"87"),
   911 => (x"a3",x"cb",x"4b",x"bf"),
   912 => (x"cf",x"4c",x"11",x"49"),
   913 => (x"d2",x"c1",x"05",x"ac"),
   914 => (x"df",x"49",x"75",x"87"),
   915 => (x"cd",x"89",x"c1",x"99"),
   916 => (x"cc",x"ef",x"c2",x"91"),
   917 => (x"4a",x"a3",x"c1",x"81"),
   918 => (x"a3",x"c3",x"51",x"12"),
   919 => (x"c5",x"51",x"12",x"4a"),
   920 => (x"51",x"12",x"4a",x"a3"),
   921 => (x"12",x"4a",x"a3",x"c7"),
   922 => (x"4a",x"a3",x"c9",x"51"),
   923 => (x"a3",x"ce",x"51",x"12"),
   924 => (x"d0",x"51",x"12",x"4a"),
   925 => (x"51",x"12",x"4a",x"a3"),
   926 => (x"12",x"4a",x"a3",x"d2"),
   927 => (x"4a",x"a3",x"d4",x"51"),
   928 => (x"a3",x"d6",x"51",x"12"),
   929 => (x"d8",x"51",x"12",x"4a"),
   930 => (x"51",x"12",x"4a",x"a3"),
   931 => (x"12",x"4a",x"a3",x"dc"),
   932 => (x"4a",x"a3",x"de",x"51"),
   933 => (x"7e",x"c1",x"51",x"12"),
   934 => (x"74",x"87",x"fc",x"c0"),
   935 => (x"05",x"99",x"c8",x"49"),
   936 => (x"74",x"87",x"ed",x"c0"),
   937 => (x"05",x"99",x"d0",x"49"),
   938 => (x"e0",x"c0",x"87",x"d3"),
   939 => (x"cc",x"c0",x"02",x"66"),
   940 => (x"c0",x"49",x"73",x"87"),
   941 => (x"70",x"0f",x"66",x"e0"),
   942 => (x"d3",x"c0",x"02",x"98"),
   943 => (x"c0",x"05",x"6e",x"87"),
   944 => (x"ef",x"c2",x"87",x"c6"),
   945 => (x"50",x"c0",x"48",x"cc"),
   946 => (x"bf",x"cc",x"fe",x"c0"),
   947 => (x"87",x"e9",x"c2",x"48"),
   948 => (x"48",x"d9",x"ef",x"c2"),
   949 => (x"c2",x"7e",x"50",x"c0"),
   950 => (x"49",x"bf",x"c8",x"ef"),
   951 => (x"bf",x"f8",x"e6",x"c2"),
   952 => (x"04",x"aa",x"71",x"4a"),
   953 => (x"cf",x"87",x"f4",x"fb"),
   954 => (x"f8",x"ff",x"ff",x"ff"),
   955 => (x"fc",x"f3",x"c2",x"4c"),
   956 => (x"c8",x"c0",x"05",x"bf"),
   957 => (x"c4",x"ef",x"c2",x"87"),
   958 => (x"fa",x"c1",x"02",x"bf"),
   959 => (x"f4",x"e6",x"c2",x"87"),
   960 => (x"c0",x"eb",x"49",x"bf"),
   961 => (x"f8",x"e6",x"c2",x"87"),
   962 => (x"48",x"a6",x"c4",x"58"),
   963 => (x"bf",x"f4",x"e6",x"c2"),
   964 => (x"c4",x"ef",x"c2",x"78"),
   965 => (x"db",x"c0",x"02",x"bf"),
   966 => (x"49",x"66",x"c4",x"87"),
   967 => (x"a9",x"74",x"99",x"74"),
   968 => (x"87",x"c8",x"c0",x"02"),
   969 => (x"c0",x"48",x"a6",x"c8"),
   970 => (x"87",x"e7",x"c0",x"78"),
   971 => (x"c1",x"48",x"a6",x"c8"),
   972 => (x"87",x"df",x"c0",x"78"),
   973 => (x"cf",x"49",x"66",x"c4"),
   974 => (x"a9",x"99",x"f8",x"ff"),
   975 => (x"87",x"c8",x"c0",x"02"),
   976 => (x"c0",x"48",x"a6",x"cc"),
   977 => (x"87",x"c5",x"c0",x"78"),
   978 => (x"c1",x"48",x"a6",x"cc"),
   979 => (x"48",x"a6",x"c8",x"78"),
   980 => (x"c8",x"78",x"66",x"cc"),
   981 => (x"de",x"c0",x"05",x"66"),
   982 => (x"49",x"66",x"c4",x"87"),
   983 => (x"ee",x"c2",x"89",x"c2"),
   984 => (x"c2",x"91",x"bf",x"fc"),
   985 => (x"48",x"bf",x"e0",x"f3"),
   986 => (x"e6",x"c2",x"80",x"71"),
   987 => (x"e6",x"c2",x"58",x"f4"),
   988 => (x"78",x"c0",x"48",x"f8"),
   989 => (x"c0",x"87",x"d4",x"f9"),
   990 => (x"ff",x"ff",x"cf",x"48"),
   991 => (x"f0",x"4c",x"f8",x"ff"),
   992 => (x"26",x"4d",x"26",x"8e"),
   993 => (x"26",x"4b",x"26",x"4c"),
   994 => (x"00",x"00",x"00",x"4f"),
   995 => (x"00",x"00",x"00",x"00"),
   996 => (x"ff",x"ff",x"ff",x"ff"),
   997 => (x"48",x"d4",x"ff",x"1e"),
   998 => (x"26",x"78",x"ff",x"c3"),
   999 => (x"d4",x"ff",x"1e",x"4f"),
  1000 => (x"78",x"ff",x"c3",x"48"),
  1001 => (x"c0",x"48",x"d0",x"ff"),
  1002 => (x"d4",x"ff",x"78",x"e1"),
  1003 => (x"26",x"78",x"d4",x"48"),
  1004 => (x"d0",x"ff",x"1e",x"4f"),
  1005 => (x"78",x"e0",x"c0",x"48"),
  1006 => (x"ff",x"1e",x"4f",x"26"),
  1007 => (x"49",x"70",x"87",x"d6"),
  1008 => (x"87",x"c6",x"02",x"99"),
  1009 => (x"05",x"a9",x"fb",x"c0"),
  1010 => (x"48",x"71",x"87",x"f1"),
  1011 => (x"5e",x"0e",x"4f",x"26"),
  1012 => (x"71",x"0e",x"5c",x"5b"),
  1013 => (x"fe",x"4c",x"c0",x"4b"),
  1014 => (x"49",x"70",x"87",x"fa"),
  1015 => (x"f9",x"c0",x"02",x"99"),
  1016 => (x"a9",x"ec",x"c0",x"87"),
  1017 => (x"87",x"f2",x"c0",x"02"),
  1018 => (x"02",x"a9",x"fb",x"c0"),
  1019 => (x"cc",x"87",x"eb",x"c0"),
  1020 => (x"03",x"ac",x"b7",x"66"),
  1021 => (x"66",x"d0",x"87",x"c7"),
  1022 => (x"71",x"87",x"c2",x"02"),
  1023 => (x"02",x"99",x"71",x"53"),
  1024 => (x"84",x"c1",x"87",x"c2"),
  1025 => (x"70",x"87",x"cd",x"fe"),
  1026 => (x"cd",x"02",x"99",x"49"),
  1027 => (x"a9",x"ec",x"c0",x"87"),
  1028 => (x"c0",x"87",x"c7",x"02"),
  1029 => (x"ff",x"05",x"a9",x"fb"),
  1030 => (x"66",x"d0",x"87",x"d5"),
  1031 => (x"c0",x"87",x"c3",x"02"),
  1032 => (x"fb",x"c0",x"7b",x"97"),
  1033 => (x"87",x"c7",x"05",x"a9"),
  1034 => (x"0a",x"c0",x"4a",x"74"),
  1035 => (x"74",x"87",x"c2",x"8a"),
  1036 => (x"26",x"48",x"72",x"4a"),
  1037 => (x"26",x"4b",x"26",x"4c"),
  1038 => (x"d7",x"fd",x"1e",x"4f"),
  1039 => (x"c0",x"49",x"70",x"87"),
  1040 => (x"c9",x"04",x"a9",x"f0"),
  1041 => (x"a9",x"f9",x"c0",x"87"),
  1042 => (x"c0",x"87",x"c3",x"01"),
  1043 => (x"c1",x"c1",x"89",x"f0"),
  1044 => (x"87",x"c9",x"04",x"a9"),
  1045 => (x"01",x"a9",x"da",x"c1"),
  1046 => (x"f7",x"c0",x"87",x"c3"),
  1047 => (x"26",x"48",x"71",x"89"),
  1048 => (x"5b",x"5e",x"0e",x"4f"),
  1049 => (x"f8",x"0e",x"5d",x"5c"),
  1050 => (x"c0",x"4c",x"71",x"86"),
  1051 => (x"87",x"ed",x"fc",x"7e"),
  1052 => (x"c4",x"c1",x"4b",x"c0"),
  1053 => (x"49",x"bf",x"97",x"c0"),
  1054 => (x"cf",x"04",x"a9",x"c0"),
  1055 => (x"87",x"fa",x"fc",x"87"),
  1056 => (x"c4",x"c1",x"83",x"c1"),
  1057 => (x"49",x"bf",x"97",x"c0"),
  1058 => (x"87",x"f1",x"06",x"ab"),
  1059 => (x"97",x"c0",x"c4",x"c1"),
  1060 => (x"87",x"cf",x"02",x"bf"),
  1061 => (x"70",x"87",x"fd",x"fb"),
  1062 => (x"c6",x"02",x"99",x"49"),
  1063 => (x"a9",x"ec",x"c0",x"87"),
  1064 => (x"c0",x"87",x"f1",x"05"),
  1065 => (x"87",x"ec",x"fb",x"4b"),
  1066 => (x"e7",x"fb",x"4d",x"70"),
  1067 => (x"58",x"a6",x"c8",x"87"),
  1068 => (x"70",x"87",x"e1",x"fb"),
  1069 => (x"c8",x"83",x"c1",x"4a"),
  1070 => (x"69",x"97",x"49",x"a4"),
  1071 => (x"da",x"05",x"ad",x"49"),
  1072 => (x"49",x"a4",x"c9",x"87"),
  1073 => (x"c4",x"49",x"69",x"97"),
  1074 => (x"ce",x"05",x"a9",x"66"),
  1075 => (x"49",x"a4",x"ca",x"87"),
  1076 => (x"aa",x"49",x"69",x"97"),
  1077 => (x"c1",x"87",x"c4",x"05"),
  1078 => (x"c0",x"87",x"d0",x"7e"),
  1079 => (x"c6",x"02",x"ad",x"ec"),
  1080 => (x"ad",x"fb",x"c0",x"87"),
  1081 => (x"c0",x"87",x"c4",x"05"),
  1082 => (x"6e",x"7e",x"c1",x"4b"),
  1083 => (x"87",x"f5",x"fe",x"02"),
  1084 => (x"73",x"87",x"fe",x"fa"),
  1085 => (x"26",x"8e",x"f8",x"48"),
  1086 => (x"26",x"4c",x"26",x"4d"),
  1087 => (x"00",x"4f",x"26",x"4b"),
  1088 => (x"1e",x"73",x"1e",x"00"),
  1089 => (x"c8",x"4b",x"d4",x"ff"),
  1090 => (x"d0",x"ff",x"4a",x"66"),
  1091 => (x"78",x"c5",x"c8",x"48"),
  1092 => (x"c1",x"48",x"d4",x"ff"),
  1093 => (x"7b",x"11",x"78",x"d4"),
  1094 => (x"f9",x"05",x"8a",x"c1"),
  1095 => (x"48",x"d0",x"ff",x"87"),
  1096 => (x"4b",x"26",x"78",x"c4"),
  1097 => (x"5e",x"0e",x"4f",x"26"),
  1098 => (x"0e",x"5d",x"5c",x"5b"),
  1099 => (x"7e",x"71",x"86",x"f8"),
  1100 => (x"f4",x"c2",x"1e",x"6e"),
  1101 => (x"c3",x"e4",x"49",x"d0"),
  1102 => (x"70",x"86",x"c4",x"87"),
  1103 => (x"ed",x"c4",x"02",x"98"),
  1104 => (x"dc",x"f1",x"c1",x"87"),
  1105 => (x"49",x"6e",x"4c",x"bf"),
  1106 => (x"c8",x"87",x"d6",x"fc"),
  1107 => (x"c9",x"c1",x"58",x"a6"),
  1108 => (x"fc",x"fe",x"1e",x"fc"),
  1109 => (x"86",x"c4",x"87",x"f6"),
  1110 => (x"87",x"c5",x"05",x"66"),
  1111 => (x"c1",x"48",x"a6",x"c4"),
  1112 => (x"48",x"d0",x"ff",x"78"),
  1113 => (x"d4",x"ff",x"78",x"c5"),
  1114 => (x"78",x"d5",x"c1",x"48"),
  1115 => (x"c1",x"49",x"66",x"c4"),
  1116 => (x"c1",x"31",x"c6",x"89"),
  1117 => (x"bf",x"97",x"d4",x"f1"),
  1118 => (x"b0",x"71",x"48",x"4a"),
  1119 => (x"78",x"08",x"d4",x"ff"),
  1120 => (x"c4",x"48",x"d0",x"ff"),
  1121 => (x"cc",x"f4",x"c2",x"78"),
  1122 => (x"d0",x"49",x"bf",x"97"),
  1123 => (x"87",x"dd",x"02",x"99"),
  1124 => (x"d4",x"ff",x"78",x"c5"),
  1125 => (x"78",x"d6",x"c1",x"48"),
  1126 => (x"d4",x"ff",x"4a",x"c0"),
  1127 => (x"78",x"ff",x"c3",x"48"),
  1128 => (x"e0",x"c0",x"82",x"c1"),
  1129 => (x"87",x"f2",x"04",x"aa"),
  1130 => (x"c4",x"48",x"d0",x"ff"),
  1131 => (x"48",x"d4",x"ff",x"78"),
  1132 => (x"ff",x"78",x"ff",x"c3"),
  1133 => (x"78",x"c5",x"48",x"d0"),
  1134 => (x"c1",x"48",x"d4",x"ff"),
  1135 => (x"78",x"c1",x"78",x"d3"),
  1136 => (x"c4",x"48",x"d0",x"ff"),
  1137 => (x"ac",x"b7",x"c0",x"78"),
  1138 => (x"87",x"cb",x"c2",x"06"),
  1139 => (x"bf",x"d8",x"f4",x"c2"),
  1140 => (x"7e",x"74",x"8c",x"4b"),
  1141 => (x"c1",x"02",x"9b",x"73"),
  1142 => (x"c0",x"c8",x"87",x"dd"),
  1143 => (x"b7",x"c0",x"8b",x"4d"),
  1144 => (x"87",x"c6",x"03",x"ab"),
  1145 => (x"4d",x"a3",x"c0",x"c8"),
  1146 => (x"f4",x"c2",x"4b",x"c0"),
  1147 => (x"49",x"bf",x"97",x"cc"),
  1148 => (x"cf",x"02",x"99",x"d0"),
  1149 => (x"c2",x"1e",x"c0",x"87"),
  1150 => (x"e5",x"49",x"d0",x"f4"),
  1151 => (x"86",x"c4",x"87",x"f2"),
  1152 => (x"87",x"d8",x"4c",x"70"),
  1153 => (x"1e",x"fc",x"e6",x"c2"),
  1154 => (x"49",x"d0",x"f4",x"c2"),
  1155 => (x"70",x"87",x"e1",x"e5"),
  1156 => (x"c2",x"1e",x"75",x"4c"),
  1157 => (x"fb",x"49",x"fc",x"e6"),
  1158 => (x"86",x"c8",x"87",x"e7"),
  1159 => (x"c5",x"05",x"9c",x"74"),
  1160 => (x"c1",x"48",x"c0",x"87"),
  1161 => (x"1e",x"c1",x"87",x"ca"),
  1162 => (x"49",x"d0",x"f4",x"c2"),
  1163 => (x"c4",x"87",x"f4",x"e3"),
  1164 => (x"05",x"9b",x"73",x"86"),
  1165 => (x"6e",x"87",x"e3",x"fe"),
  1166 => (x"ac",x"b7",x"c0",x"4c"),
  1167 => (x"c2",x"87",x"d1",x"06"),
  1168 => (x"c0",x"48",x"d0",x"f4"),
  1169 => (x"c0",x"80",x"d0",x"78"),
  1170 => (x"c2",x"80",x"f4",x"78"),
  1171 => (x"78",x"bf",x"dc",x"f4"),
  1172 => (x"01",x"ac",x"b7",x"c0"),
  1173 => (x"ff",x"87",x"f5",x"fd"),
  1174 => (x"78",x"c5",x"48",x"d0"),
  1175 => (x"c1",x"48",x"d4",x"ff"),
  1176 => (x"78",x"c0",x"78",x"d3"),
  1177 => (x"c4",x"48",x"d0",x"ff"),
  1178 => (x"c0",x"48",x"c1",x"78"),
  1179 => (x"48",x"c0",x"87",x"c2"),
  1180 => (x"4d",x"26",x"8e",x"f8"),
  1181 => (x"4b",x"26",x"4c",x"26"),
  1182 => (x"00",x"00",x"4f",x"26"),
  1183 => (x"20",x"74",x"6f",x"47"),
  1184 => (x"69",x"74",x"78",x"65"),
  1185 => (x"00",x"00",x"64",x"6e"),
  1186 => (x"64",x"61",x"6f",x"4c"),
  1187 => (x"2e",x"67",x"6e",x"69"),
  1188 => (x"00",x"00",x"2e",x"2e"),
  1189 => (x"61",x"42",x"20",x"80"),
  1190 => (x"00",x"00",x"6b",x"63"),
  1191 => (x"64",x"61",x"6f",x"4c"),
  1192 => (x"20",x"2e",x"2a",x"20"),
  1193 => (x"00",x"00",x"00",x"00"),
  1194 => (x"00",x"00",x"20",x"3a"),
  1195 => (x"61",x"42",x"20",x"80"),
  1196 => (x"00",x"00",x"6b",x"63"),
  1197 => (x"78",x"45",x"20",x"80"),
  1198 => (x"00",x"00",x"74",x"69"),
  1199 => (x"49",x"20",x"44",x"53"),
  1200 => (x"2e",x"74",x"69",x"6e"),
  1201 => (x"00",x"00",x"00",x"2e"),
  1202 => (x"00",x"00",x"4b",x"4f"),
  1203 => (x"54",x"4f",x"4f",x"42"),
  1204 => (x"20",x"20",x"20",x"20"),
  1205 => (x"00",x"4d",x"4f",x"52"),
  1206 => (x"5c",x"5b",x"5e",x"0e"),
  1207 => (x"86",x"fc",x"0e",x"5d"),
  1208 => (x"4b",x"c0",x"4d",x"71"),
  1209 => (x"c0",x"04",x"ad",x"4c"),
  1210 => (x"c1",x"c1",x"87",x"e8"),
  1211 => (x"9c",x"74",x"1e",x"e1"),
  1212 => (x"c0",x"87",x"c4",x"02"),
  1213 => (x"c1",x"87",x"c2",x"4a"),
  1214 => (x"ea",x"49",x"72",x"4a"),
  1215 => (x"86",x"c4",x"87",x"d7"),
  1216 => (x"83",x"c1",x"7e",x"70"),
  1217 => (x"87",x"c2",x"05",x"6e"),
  1218 => (x"84",x"c1",x"4b",x"75"),
  1219 => (x"ff",x"06",x"ab",x"75"),
  1220 => (x"48",x"6e",x"87",x"d8"),
  1221 => (x"4d",x"26",x"8e",x"fc"),
  1222 => (x"4b",x"26",x"4c",x"26"),
  1223 => (x"5e",x"0e",x"4f",x"26"),
  1224 => (x"0e",x"5d",x"5c",x"5b"),
  1225 => (x"4d",x"71",x"86",x"f4"),
  1226 => (x"c2",x"91",x"de",x"49"),
  1227 => (x"71",x"48",x"f0",x"f5"),
  1228 => (x"6e",x"7e",x"70",x"80"),
  1229 => (x"c2",x"02",x"bf",x"97"),
  1230 => (x"f5",x"c2",x"87",x"cb"),
  1231 => (x"75",x"49",x"bf",x"e0"),
  1232 => (x"d3",x"fe",x"71",x"81"),
  1233 => (x"58",x"a6",x"c8",x"87"),
  1234 => (x"c1",x"02",x"66",x"c4"),
  1235 => (x"f5",x"c2",x"87",x"e1"),
  1236 => (x"66",x"c4",x"4b",x"e4"),
  1237 => (x"fe",x"49",x"cb",x"4a"),
  1238 => (x"75",x"87",x"c7",x"fb"),
  1239 => (x"c1",x"93",x"cc",x"4b"),
  1240 => (x"c4",x"83",x"e0",x"f1"),
  1241 => (x"c8",x"ca",x"c1",x"83"),
  1242 => (x"c1",x"49",x"75",x"7b"),
  1243 => (x"6e",x"87",x"fd",x"c0"),
  1244 => (x"d8",x"f1",x"c1",x"7b"),
  1245 => (x"cc",x"48",x"bf",x"97"),
  1246 => (x"98",x"70",x"58",x"a6"),
  1247 => (x"48",x"87",x"db",x"02"),
  1248 => (x"70",x"88",x"f0",x"c0"),
  1249 => (x"02",x"98",x"48",x"7e"),
  1250 => (x"c1",x"4c",x"87",x"d9"),
  1251 => (x"87",x"d3",x"02",x"8c"),
  1252 => (x"87",x"cf",x"02",x"8c"),
  1253 => (x"87",x"cb",x"02",x"8c"),
  1254 => (x"f5",x"c2",x"87",x"d5"),
  1255 => (x"c5",x"f6",x"49",x"e4"),
  1256 => (x"6e",x"87",x"cc",x"87"),
  1257 => (x"e4",x"f5",x"c2",x"1e"),
  1258 => (x"f3",x"d4",x"c1",x"49"),
  1259 => (x"75",x"86",x"c4",x"87"),
  1260 => (x"f7",x"ff",x"c0",x"49"),
  1261 => (x"c1",x"49",x"c0",x"87"),
  1262 => (x"c2",x"87",x"d2",x"c1"),
  1263 => (x"c0",x"48",x"c8",x"f4"),
  1264 => (x"e2",x"df",x"49",x"50"),
  1265 => (x"26",x"8e",x"f4",x"87"),
  1266 => (x"26",x"4c",x"26",x"4d"),
  1267 => (x"1e",x"4f",x"26",x"4b"),
  1268 => (x"4b",x"71",x"1e",x"73"),
  1269 => (x"e0",x"f5",x"c2",x"49"),
  1270 => (x"fb",x"71",x"81",x"bf"),
  1271 => (x"4a",x"70",x"87",x"fa"),
  1272 => (x"87",x"c4",x"02",x"9a"),
  1273 => (x"87",x"e7",x"e4",x"49"),
  1274 => (x"48",x"e0",x"f5",x"c2"),
  1275 => (x"49",x"73",x"78",x"c0"),
  1276 => (x"26",x"87",x"fa",x"c1"),
  1277 => (x"1e",x"4f",x"26",x"4b"),
  1278 => (x"4b",x"71",x"1e",x"73"),
  1279 => (x"02",x"4a",x"a3",x"c4"),
  1280 => (x"c1",x"87",x"d0",x"c1"),
  1281 => (x"87",x"dc",x"02",x"8a"),
  1282 => (x"f2",x"c0",x"02",x"8a"),
  1283 => (x"c1",x"05",x"8a",x"87"),
  1284 => (x"f5",x"c2",x"87",x"d3"),
  1285 => (x"c1",x"02",x"bf",x"e0"),
  1286 => (x"c1",x"48",x"87",x"cb"),
  1287 => (x"e4",x"f5",x"c2",x"88"),
  1288 => (x"87",x"c1",x"c1",x"58"),
  1289 => (x"bf",x"e0",x"f5",x"c2"),
  1290 => (x"c2",x"89",x"c6",x"49"),
  1291 => (x"c0",x"59",x"e4",x"f5"),
  1292 => (x"c0",x"03",x"a9",x"b7"),
  1293 => (x"f5",x"c2",x"87",x"ef"),
  1294 => (x"78",x"c0",x"48",x"e0"),
  1295 => (x"c2",x"87",x"e6",x"c0"),
  1296 => (x"02",x"bf",x"dc",x"f5"),
  1297 => (x"f5",x"c2",x"87",x"df"),
  1298 => (x"c1",x"48",x"bf",x"e0"),
  1299 => (x"e4",x"f5",x"c2",x"80"),
  1300 => (x"c2",x"87",x"d2",x"58"),
  1301 => (x"02",x"bf",x"dc",x"f5"),
  1302 => (x"f5",x"c2",x"87",x"cb"),
  1303 => (x"c6",x"48",x"bf",x"e0"),
  1304 => (x"e4",x"f5",x"c2",x"80"),
  1305 => (x"c4",x"49",x"73",x"58"),
  1306 => (x"26",x"4b",x"26",x"87"),
  1307 => (x"5b",x"5e",x"0e",x"4f"),
  1308 => (x"f0",x"0e",x"5d",x"5c"),
  1309 => (x"59",x"a6",x"d0",x"86"),
  1310 => (x"4d",x"fc",x"e6",x"c2"),
  1311 => (x"f5",x"c2",x"4c",x"c0"),
  1312 => (x"78",x"c1",x"48",x"dc"),
  1313 => (x"c0",x"48",x"a6",x"c8"),
  1314 => (x"c2",x"7e",x"75",x"78"),
  1315 => (x"48",x"bf",x"e0",x"f5"),
  1316 => (x"c1",x"06",x"a8",x"c0"),
  1317 => (x"a6",x"c8",x"87",x"c0"),
  1318 => (x"c2",x"7e",x"75",x"5c"),
  1319 => (x"98",x"48",x"fc",x"e6"),
  1320 => (x"87",x"f2",x"c0",x"02"),
  1321 => (x"c1",x"4d",x"66",x"c4"),
  1322 => (x"cc",x"1e",x"e1",x"c1"),
  1323 => (x"87",x"c4",x"02",x"66"),
  1324 => (x"87",x"c2",x"4c",x"c0"),
  1325 => (x"49",x"74",x"4c",x"c1"),
  1326 => (x"c4",x"87",x"da",x"e3"),
  1327 => (x"c1",x"7e",x"70",x"86"),
  1328 => (x"48",x"66",x"c8",x"85"),
  1329 => (x"a6",x"cc",x"80",x"c1"),
  1330 => (x"e0",x"f5",x"c2",x"58"),
  1331 => (x"c5",x"03",x"ad",x"bf"),
  1332 => (x"ff",x"05",x"6e",x"87"),
  1333 => (x"4d",x"6e",x"87",x"d1"),
  1334 => (x"9d",x"75",x"4c",x"c0"),
  1335 => (x"87",x"dc",x"c3",x"02"),
  1336 => (x"1e",x"e1",x"c1",x"c1"),
  1337 => (x"c7",x"02",x"66",x"cc"),
  1338 => (x"48",x"a6",x"c8",x"87"),
  1339 => (x"87",x"c5",x"78",x"c0"),
  1340 => (x"c1",x"48",x"a6",x"c8"),
  1341 => (x"49",x"66",x"c8",x"78"),
  1342 => (x"c4",x"87",x"da",x"e2"),
  1343 => (x"48",x"7e",x"70",x"86"),
  1344 => (x"e4",x"c2",x"02",x"98"),
  1345 => (x"81",x"cb",x"49",x"87"),
  1346 => (x"d0",x"49",x"69",x"97"),
  1347 => (x"d4",x"c1",x"02",x"99"),
  1348 => (x"cc",x"49",x"74",x"87"),
  1349 => (x"e0",x"f1",x"c1",x"91"),
  1350 => (x"cf",x"cf",x"c1",x"81"),
  1351 => (x"c3",x"81",x"c8",x"79"),
  1352 => (x"49",x"74",x"51",x"ff"),
  1353 => (x"f5",x"c2",x"91",x"de"),
  1354 => (x"85",x"71",x"4d",x"f0"),
  1355 => (x"7d",x"97",x"c1",x"c2"),
  1356 => (x"c0",x"49",x"a5",x"c1"),
  1357 => (x"ef",x"c2",x"51",x"e0"),
  1358 => (x"02",x"bf",x"97",x"cc"),
  1359 => (x"84",x"c1",x"87",x"d2"),
  1360 => (x"c2",x"4b",x"a5",x"c2"),
  1361 => (x"db",x"4a",x"cc",x"ef"),
  1362 => (x"d5",x"f3",x"fe",x"49"),
  1363 => (x"87",x"d9",x"c1",x"87"),
  1364 => (x"c0",x"49",x"a5",x"cd"),
  1365 => (x"c2",x"84",x"c1",x"51"),
  1366 => (x"4a",x"6e",x"4b",x"a5"),
  1367 => (x"f3",x"fe",x"49",x"cb"),
  1368 => (x"c4",x"c1",x"87",x"c0"),
  1369 => (x"cc",x"49",x"74",x"87"),
  1370 => (x"e0",x"f1",x"c1",x"91"),
  1371 => (x"de",x"cc",x"c1",x"81"),
  1372 => (x"cc",x"ef",x"c2",x"79"),
  1373 => (x"d8",x"02",x"bf",x"97"),
  1374 => (x"de",x"49",x"74",x"87"),
  1375 => (x"c2",x"84",x"c1",x"91"),
  1376 => (x"71",x"4b",x"f0",x"f5"),
  1377 => (x"cc",x"ef",x"c2",x"83"),
  1378 => (x"fe",x"49",x"dd",x"4a"),
  1379 => (x"d8",x"87",x"d3",x"f2"),
  1380 => (x"de",x"4b",x"74",x"87"),
  1381 => (x"f0",x"f5",x"c2",x"93"),
  1382 => (x"49",x"a3",x"cb",x"83"),
  1383 => (x"84",x"c1",x"51",x"c0"),
  1384 => (x"cb",x"4a",x"6e",x"73"),
  1385 => (x"f9",x"f1",x"fe",x"49"),
  1386 => (x"48",x"66",x"c8",x"87"),
  1387 => (x"a6",x"cc",x"80",x"c1"),
  1388 => (x"03",x"ac",x"c7",x"58"),
  1389 => (x"6e",x"87",x"c5",x"c0"),
  1390 => (x"87",x"e4",x"fc",x"05"),
  1391 => (x"c0",x"03",x"ac",x"c7"),
  1392 => (x"f5",x"c2",x"87",x"e4"),
  1393 => (x"78",x"c0",x"48",x"dc"),
  1394 => (x"91",x"cc",x"49",x"74"),
  1395 => (x"81",x"e0",x"f1",x"c1"),
  1396 => (x"79",x"de",x"cc",x"c1"),
  1397 => (x"91",x"de",x"49",x"74"),
  1398 => (x"81",x"f0",x"f5",x"c2"),
  1399 => (x"84",x"c1",x"51",x"c0"),
  1400 => (x"ff",x"04",x"ac",x"c7"),
  1401 => (x"f2",x"c1",x"87",x"dc"),
  1402 => (x"50",x"c0",x"48",x"fc"),
  1403 => (x"d9",x"c1",x"80",x"f7"),
  1404 => (x"ca",x"c1",x"40",x"c5"),
  1405 => (x"80",x"c8",x"78",x"d4"),
  1406 => (x"78",x"f7",x"cf",x"c1"),
  1407 => (x"c0",x"49",x"66",x"cc"),
  1408 => (x"f0",x"87",x"e9",x"f6"),
  1409 => (x"26",x"4d",x"26",x"8e"),
  1410 => (x"26",x"4b",x"26",x"4c"),
  1411 => (x"1e",x"73",x"1e",x"4f"),
  1412 => (x"cc",x"49",x"4b",x"71"),
  1413 => (x"e0",x"f1",x"c1",x"91"),
  1414 => (x"4a",x"a1",x"c8",x"81"),
  1415 => (x"48",x"d4",x"f1",x"c1"),
  1416 => (x"a1",x"c9",x"50",x"12"),
  1417 => (x"c0",x"c4",x"c1",x"4a"),
  1418 => (x"ca",x"50",x"12",x"48"),
  1419 => (x"d8",x"f1",x"c1",x"81"),
  1420 => (x"73",x"50",x"11",x"48"),
  1421 => (x"87",x"f5",x"f8",x"49"),
  1422 => (x"4f",x"26",x"4b",x"26"),
  1423 => (x"c0",x"49",x"c0",x"1e"),
  1424 => (x"26",x"87",x"ca",x"f7"),
  1425 => (x"4a",x"71",x"1e",x"4f"),
  1426 => (x"c1",x"91",x"cc",x"49"),
  1427 => (x"c8",x"81",x"e0",x"f1"),
  1428 => (x"c8",x"f4",x"c2",x"81"),
  1429 => (x"c0",x"50",x"11",x"48"),
  1430 => (x"fe",x"49",x"a2",x"f0"),
  1431 => (x"c0",x"87",x"cf",x"ed"),
  1432 => (x"87",x"c3",x"d5",x"49"),
  1433 => (x"ff",x"1e",x"4f",x"26"),
  1434 => (x"ff",x"c3",x"4a",x"d4"),
  1435 => (x"48",x"d0",x"ff",x"7a"),
  1436 => (x"de",x"78",x"e1",x"c0"),
  1437 => (x"48",x"7a",x"71",x"7a"),
  1438 => (x"70",x"28",x"b7",x"c8"),
  1439 => (x"d0",x"48",x"71",x"7a"),
  1440 => (x"7a",x"70",x"28",x"b7"),
  1441 => (x"b7",x"d8",x"48",x"71"),
  1442 => (x"ff",x"7a",x"70",x"28"),
  1443 => (x"e0",x"c0",x"48",x"d0"),
  1444 => (x"0e",x"4f",x"26",x"78"),
  1445 => (x"5d",x"5c",x"5b",x"5e"),
  1446 => (x"71",x"86",x"f4",x"0e"),
  1447 => (x"91",x"cc",x"49",x"4d"),
  1448 => (x"81",x"e0",x"f1",x"c1"),
  1449 => (x"ca",x"4a",x"a1",x"c8"),
  1450 => (x"a6",x"c4",x"7e",x"a1"),
  1451 => (x"c4",x"f4",x"c2",x"48"),
  1452 => (x"97",x"6e",x"78",x"bf"),
  1453 => (x"66",x"c4",x"4b",x"bf"),
  1454 => (x"12",x"2c",x"73",x"4c"),
  1455 => (x"58",x"a6",x"cc",x"48"),
  1456 => (x"84",x"c1",x"9c",x"70"),
  1457 => (x"69",x"97",x"81",x"c9"),
  1458 => (x"04",x"ac",x"b7",x"49"),
  1459 => (x"4c",x"c0",x"87",x"c2"),
  1460 => (x"4a",x"bf",x"97",x"6e"),
  1461 => (x"72",x"49",x"66",x"c8"),
  1462 => (x"c4",x"b9",x"ff",x"31"),
  1463 => (x"48",x"74",x"99",x"66"),
  1464 => (x"4a",x"70",x"30",x"72"),
  1465 => (x"c8",x"f4",x"c2",x"b1"),
  1466 => (x"f9",x"fd",x"71",x"59"),
  1467 => (x"c2",x"1e",x"c7",x"87"),
  1468 => (x"1e",x"bf",x"d8",x"f5"),
  1469 => (x"1e",x"e0",x"f1",x"c1"),
  1470 => (x"97",x"c8",x"f4",x"c2"),
  1471 => (x"f4",x"c1",x"49",x"bf"),
  1472 => (x"c0",x"49",x"75",x"87"),
  1473 => (x"e8",x"87",x"e5",x"f2"),
  1474 => (x"26",x"4d",x"26",x"8e"),
  1475 => (x"26",x"4b",x"26",x"4c"),
  1476 => (x"1e",x"73",x"1e",x"4f"),
  1477 => (x"fd",x"49",x"4b",x"71"),
  1478 => (x"49",x"73",x"87",x"f9"),
  1479 => (x"26",x"87",x"f4",x"fd"),
  1480 => (x"1e",x"4f",x"26",x"4b"),
  1481 => (x"4b",x"71",x"1e",x"73"),
  1482 => (x"02",x"4a",x"a3",x"c2"),
  1483 => (x"8a",x"c1",x"87",x"d6"),
  1484 => (x"87",x"e2",x"c0",x"05"),
  1485 => (x"bf",x"d8",x"f5",x"c2"),
  1486 => (x"48",x"87",x"db",x"02"),
  1487 => (x"f5",x"c2",x"88",x"c1"),
  1488 => (x"87",x"d2",x"58",x"dc"),
  1489 => (x"bf",x"dc",x"f5",x"c2"),
  1490 => (x"c2",x"87",x"cb",x"02"),
  1491 => (x"48",x"bf",x"d8",x"f5"),
  1492 => (x"f5",x"c2",x"80",x"c1"),
  1493 => (x"1e",x"c7",x"58",x"dc"),
  1494 => (x"bf",x"d8",x"f5",x"c2"),
  1495 => (x"e0",x"f1",x"c1",x"1e"),
  1496 => (x"c8",x"f4",x"c2",x"1e"),
  1497 => (x"cc",x"49",x"bf",x"97"),
  1498 => (x"c0",x"49",x"73",x"87"),
  1499 => (x"f4",x"87",x"fd",x"f0"),
  1500 => (x"26",x"4b",x"26",x"8e"),
  1501 => (x"5b",x"5e",x"0e",x"4f"),
  1502 => (x"ff",x"0e",x"5d",x"5c"),
  1503 => (x"e8",x"c0",x"86",x"cc"),
  1504 => (x"a6",x"cc",x"59",x"a6"),
  1505 => (x"c4",x"78",x"c0",x"48"),
  1506 => (x"c4",x"78",x"c0",x"80"),
  1507 => (x"c4",x"78",x"c0",x"80"),
  1508 => (x"66",x"c8",x"c1",x"80"),
  1509 => (x"c1",x"80",x"c4",x"78"),
  1510 => (x"c1",x"80",x"c4",x"78"),
  1511 => (x"dc",x"f5",x"c2",x"78"),
  1512 => (x"ff",x"78",x"c1",x"48"),
  1513 => (x"e0",x"87",x"f6",x"df"),
  1514 => (x"df",x"ff",x"87",x"d0"),
  1515 => (x"4d",x"70",x"87",x"e6"),
  1516 => (x"02",x"ad",x"fb",x"c0"),
  1517 => (x"c0",x"87",x"f3",x"c1"),
  1518 => (x"c1",x"05",x"66",x"e4"),
  1519 => (x"c4",x"c1",x"87",x"e8"),
  1520 => (x"82",x"c4",x"4a",x"66"),
  1521 => (x"ca",x"c1",x"7e",x"6a"),
  1522 => (x"49",x"6e",x"48",x"dc"),
  1523 => (x"41",x"20",x"41",x"20"),
  1524 => (x"c4",x"c1",x"51",x"10"),
  1525 => (x"d8",x"c1",x"48",x"66"),
  1526 => (x"49",x"6a",x"78",x"cd"),
  1527 => (x"51",x"75",x"81",x"c7"),
  1528 => (x"49",x"66",x"c4",x"c1"),
  1529 => (x"51",x"c1",x"81",x"c8"),
  1530 => (x"c2",x"48",x"a6",x"dc"),
  1531 => (x"66",x"c4",x"c1",x"78"),
  1532 => (x"c0",x"81",x"c9",x"49"),
  1533 => (x"66",x"c4",x"c1",x"51"),
  1534 => (x"c0",x"81",x"ca",x"49"),
  1535 => (x"d8",x"1e",x"c1",x"51"),
  1536 => (x"c8",x"49",x"6a",x"1e"),
  1537 => (x"c5",x"df",x"ff",x"81"),
  1538 => (x"c1",x"86",x"c8",x"87"),
  1539 => (x"c0",x"48",x"66",x"c8"),
  1540 => (x"87",x"c7",x"01",x"a8"),
  1541 => (x"c1",x"48",x"a6",x"d4"),
  1542 => (x"c1",x"87",x"cf",x"78"),
  1543 => (x"c1",x"48",x"66",x"c8"),
  1544 => (x"58",x"a6",x"dc",x"88"),
  1545 => (x"de",x"ff",x"87",x"c4"),
  1546 => (x"9d",x"75",x"87",x"d0"),
  1547 => (x"87",x"f1",x"cb",x"02"),
  1548 => (x"c1",x"48",x"66",x"d4"),
  1549 => (x"03",x"a8",x"66",x"cc"),
  1550 => (x"c0",x"87",x"e6",x"cb"),
  1551 => (x"d3",x"dd",x"ff",x"7e"),
  1552 => (x"48",x"4d",x"70",x"87"),
  1553 => (x"c8",x"88",x"c6",x"c1"),
  1554 => (x"98",x"70",x"58",x"a6"),
  1555 => (x"87",x"d6",x"c1",x"02"),
  1556 => (x"c8",x"88",x"c9",x"48"),
  1557 => (x"98",x"70",x"58",x"a6"),
  1558 => (x"87",x"d7",x"c5",x"02"),
  1559 => (x"c8",x"88",x"c1",x"48"),
  1560 => (x"98",x"70",x"58",x"a6"),
  1561 => (x"87",x"f8",x"c2",x"02"),
  1562 => (x"c8",x"88",x"c3",x"48"),
  1563 => (x"98",x"70",x"58",x"a6"),
  1564 => (x"48",x"87",x"cf",x"02"),
  1565 => (x"a6",x"c8",x"88",x"c1"),
  1566 => (x"02",x"98",x"70",x"58"),
  1567 => (x"c9",x"87",x"f4",x"c4"),
  1568 => (x"f0",x"c0",x"87",x"fe"),
  1569 => (x"cb",x"dc",x"ff",x"7e"),
  1570 => (x"c0",x"4d",x"70",x"87"),
  1571 => (x"c2",x"02",x"ad",x"ec"),
  1572 => (x"c0",x"7e",x"75",x"87"),
  1573 => (x"cd",x"02",x"ad",x"ec"),
  1574 => (x"f7",x"db",x"ff",x"87"),
  1575 => (x"c0",x"4d",x"70",x"87"),
  1576 => (x"ff",x"05",x"ad",x"ec"),
  1577 => (x"e4",x"c0",x"87",x"f3"),
  1578 => (x"ea",x"c1",x"05",x"66"),
  1579 => (x"ad",x"ec",x"c0",x"87"),
  1580 => (x"ff",x"87",x"c4",x"02"),
  1581 => (x"c0",x"87",x"dd",x"db"),
  1582 => (x"dc",x"1e",x"ca",x"1e"),
  1583 => (x"93",x"cc",x"4b",x"66"),
  1584 => (x"83",x"66",x"cc",x"c1"),
  1585 => (x"6c",x"4c",x"a3",x"c4"),
  1586 => (x"c1",x"dc",x"ff",x"49"),
  1587 => (x"de",x"1e",x"c1",x"87"),
  1588 => (x"ff",x"49",x"6c",x"1e"),
  1589 => (x"d0",x"87",x"f7",x"db"),
  1590 => (x"cd",x"d8",x"c1",x"86"),
  1591 => (x"49",x"a3",x"c8",x"7b"),
  1592 => (x"c9",x"51",x"66",x"dc"),
  1593 => (x"e0",x"c0",x"49",x"a3"),
  1594 => (x"a3",x"ca",x"51",x"66"),
  1595 => (x"dc",x"51",x"6e",x"49"),
  1596 => (x"80",x"c1",x"48",x"66"),
  1597 => (x"58",x"a6",x"e0",x"c0"),
  1598 => (x"d8",x"48",x"66",x"d4"),
  1599 => (x"cb",x"04",x"a8",x"66"),
  1600 => (x"48",x"66",x"d4",x"87"),
  1601 => (x"a6",x"d8",x"80",x"c1"),
  1602 => (x"87",x"fa",x"c7",x"58"),
  1603 => (x"c1",x"48",x"66",x"d8"),
  1604 => (x"58",x"a6",x"dc",x"88"),
  1605 => (x"ff",x"87",x"ef",x"c7"),
  1606 => (x"70",x"87",x"df",x"da"),
  1607 => (x"87",x"e6",x"c7",x"4d"),
  1608 => (x"87",x"d5",x"dc",x"ff"),
  1609 => (x"d0",x"58",x"a6",x"d0"),
  1610 => (x"c6",x"06",x"a8",x"66"),
  1611 => (x"48",x"a6",x"d0",x"87"),
  1612 => (x"ff",x"78",x"66",x"cc"),
  1613 => (x"c0",x"87",x"c2",x"dc"),
  1614 => (x"c1",x"05",x"a8",x"ec"),
  1615 => (x"e4",x"c0",x"87",x"f5"),
  1616 => (x"e5",x"c1",x"05",x"66"),
  1617 => (x"49",x"66",x"d4",x"87"),
  1618 => (x"c4",x"c1",x"91",x"cc"),
  1619 => (x"a1",x"c4",x"81",x"66"),
  1620 => (x"c8",x"4c",x"6a",x"4a"),
  1621 => (x"66",x"cc",x"4a",x"a1"),
  1622 => (x"c5",x"d9",x"c1",x"52"),
  1623 => (x"f3",x"d8",x"ff",x"79"),
  1624 => (x"9d",x"4d",x"70",x"87"),
  1625 => (x"c0",x"87",x"da",x"02"),
  1626 => (x"d4",x"02",x"ad",x"fb"),
  1627 => (x"ff",x"54",x"75",x"87"),
  1628 => (x"70",x"87",x"e1",x"d8"),
  1629 => (x"c0",x"02",x"9d",x"4d"),
  1630 => (x"fb",x"c0",x"87",x"c7"),
  1631 => (x"ec",x"ff",x"05",x"ad"),
  1632 => (x"54",x"e0",x"c0",x"87"),
  1633 => (x"c0",x"54",x"c1",x"c2"),
  1634 => (x"66",x"d4",x"7c",x"97"),
  1635 => (x"a8",x"66",x"d8",x"48"),
  1636 => (x"87",x"cb",x"c0",x"04"),
  1637 => (x"c1",x"48",x"66",x"d4"),
  1638 => (x"58",x"a6",x"d8",x"80"),
  1639 => (x"d8",x"87",x"e7",x"c5"),
  1640 => (x"88",x"c1",x"48",x"66"),
  1641 => (x"c5",x"58",x"a6",x"dc"),
  1642 => (x"d8",x"ff",x"87",x"dc"),
  1643 => (x"4d",x"70",x"87",x"cc"),
  1644 => (x"cc",x"87",x"d3",x"c5"),
  1645 => (x"e4",x"c0",x"48",x"66"),
  1646 => (x"c4",x"05",x"a8",x"66"),
  1647 => (x"e8",x"c0",x"87",x"f4"),
  1648 => (x"78",x"c0",x"48",x"a6"),
  1649 => (x"87",x"f1",x"d9",x"ff"),
  1650 => (x"d9",x"ff",x"7e",x"70"),
  1651 => (x"f0",x"c0",x"87",x"eb"),
  1652 => (x"ec",x"c0",x"58",x"a6"),
  1653 => (x"c7",x"c0",x"05",x"a8"),
  1654 => (x"6e",x"48",x"a6",x"87"),
  1655 => (x"87",x"c4",x"c0",x"78"),
  1656 => (x"87",x"f0",x"d6",x"ff"),
  1657 => (x"cc",x"49",x"66",x"d4"),
  1658 => (x"66",x"c4",x"c1",x"91"),
  1659 => (x"c8",x"80",x"71",x"48"),
  1660 => (x"66",x"c4",x"58",x"a6"),
  1661 => (x"c4",x"82",x"c8",x"4a"),
  1662 => (x"81",x"ca",x"49",x"66"),
  1663 => (x"ec",x"c0",x"51",x"6e"),
  1664 => (x"81",x"c1",x"49",x"66"),
  1665 => (x"48",x"c1",x"89",x"6e"),
  1666 => (x"49",x"70",x"30",x"71"),
  1667 => (x"97",x"71",x"89",x"c1"),
  1668 => (x"c4",x"f4",x"c2",x"7a"),
  1669 => (x"29",x"6e",x"49",x"bf"),
  1670 => (x"48",x"4a",x"6a",x"97"),
  1671 => (x"f4",x"c0",x"98",x"71"),
  1672 => (x"66",x"c4",x"58",x"a6"),
  1673 => (x"cc",x"80",x"c4",x"48"),
  1674 => (x"66",x"c8",x"58",x"a6"),
  1675 => (x"e4",x"c0",x"4c",x"bf"),
  1676 => (x"66",x"cc",x"48",x"66"),
  1677 => (x"c5",x"c0",x"02",x"a8"),
  1678 => (x"c0",x"7e",x"c0",x"87"),
  1679 => (x"7e",x"c1",x"87",x"c2"),
  1680 => (x"e0",x"c0",x"1e",x"6e"),
  1681 => (x"ff",x"49",x"74",x"1e"),
  1682 => (x"c8",x"87",x"c3",x"d6"),
  1683 => (x"c0",x"4d",x"70",x"86"),
  1684 => (x"c1",x"06",x"ad",x"b7"),
  1685 => (x"84",x"75",x"87",x"d4"),
  1686 => (x"49",x"bf",x"66",x"c8"),
  1687 => (x"74",x"81",x"e0",x"c0"),
  1688 => (x"ca",x"c1",x"4b",x"89"),
  1689 => (x"fe",x"71",x"4a",x"e8"),
  1690 => (x"c2",x"87",x"f7",x"de"),
  1691 => (x"c0",x"7e",x"74",x"84"),
  1692 => (x"c1",x"48",x"66",x"e8"),
  1693 => (x"a6",x"ec",x"c0",x"80"),
  1694 => (x"66",x"f0",x"c0",x"58"),
  1695 => (x"70",x"81",x"c1",x"49"),
  1696 => (x"c5",x"c0",x"02",x"a9"),
  1697 => (x"c0",x"4c",x"c0",x"87"),
  1698 => (x"4c",x"c1",x"87",x"c2"),
  1699 => (x"66",x"cc",x"1e",x"74"),
  1700 => (x"e0",x"c0",x"49",x"bf"),
  1701 => (x"89",x"66",x"c4",x"81"),
  1702 => (x"66",x"c8",x"1e",x"71"),
  1703 => (x"ed",x"d4",x"ff",x"49"),
  1704 => (x"c0",x"86",x"c8",x"87"),
  1705 => (x"ff",x"01",x"a8",x"b7"),
  1706 => (x"e8",x"c0",x"87",x"c5"),
  1707 => (x"d3",x"c0",x"02",x"66"),
  1708 => (x"49",x"66",x"c4",x"87"),
  1709 => (x"e8",x"c0",x"81",x"c9"),
  1710 => (x"66",x"c4",x"51",x"66"),
  1711 => (x"d3",x"da",x"c1",x"48"),
  1712 => (x"87",x"ce",x"c0",x"78"),
  1713 => (x"c9",x"49",x"66",x"c4"),
  1714 => (x"c4",x"51",x"c2",x"81"),
  1715 => (x"dc",x"c1",x"48",x"66"),
  1716 => (x"66",x"d4",x"78",x"d1"),
  1717 => (x"a8",x"66",x"d8",x"48"),
  1718 => (x"87",x"cb",x"c0",x"04"),
  1719 => (x"c1",x"48",x"66",x"d4"),
  1720 => (x"58",x"a6",x"d8",x"80"),
  1721 => (x"d8",x"87",x"d1",x"c0"),
  1722 => (x"88",x"c1",x"48",x"66"),
  1723 => (x"c0",x"58",x"a6",x"dc"),
  1724 => (x"d3",x"ff",x"87",x"c6"),
  1725 => (x"4d",x"70",x"87",x"c4"),
  1726 => (x"c0",x"48",x"a6",x"cc"),
  1727 => (x"87",x"c6",x"c0",x"78"),
  1728 => (x"87",x"f6",x"d2",x"ff"),
  1729 => (x"e0",x"c0",x"4d",x"70"),
  1730 => (x"80",x"c1",x"48",x"66"),
  1731 => (x"58",x"a6",x"e4",x"c0"),
  1732 => (x"c0",x"02",x"9d",x"75"),
  1733 => (x"66",x"d4",x"87",x"cb"),
  1734 => (x"66",x"cc",x"c1",x"48"),
  1735 => (x"da",x"f4",x"04",x"a8"),
  1736 => (x"48",x"66",x"d4",x"87"),
  1737 => (x"c0",x"03",x"a8",x"c7"),
  1738 => (x"66",x"d4",x"87",x"e1"),
  1739 => (x"dc",x"f5",x"c2",x"4c"),
  1740 => (x"74",x"78",x"c0",x"48"),
  1741 => (x"c1",x"91",x"cc",x"49"),
  1742 => (x"c4",x"81",x"66",x"c4"),
  1743 => (x"4a",x"6a",x"4a",x"a1"),
  1744 => (x"c1",x"79",x"52",x"c0"),
  1745 => (x"04",x"ac",x"c7",x"84"),
  1746 => (x"c0",x"87",x"e2",x"ff"),
  1747 => (x"c0",x"02",x"66",x"e4"),
  1748 => (x"c4",x"c1",x"87",x"e2"),
  1749 => (x"d4",x"c1",x"49",x"66"),
  1750 => (x"66",x"c4",x"c1",x"81"),
  1751 => (x"82",x"dc",x"c1",x"4a"),
  1752 => (x"d9",x"c1",x"52",x"c0"),
  1753 => (x"c4",x"c1",x"79",x"c5"),
  1754 => (x"d8",x"c1",x"49",x"66"),
  1755 => (x"ec",x"ca",x"c1",x"81"),
  1756 => (x"87",x"d6",x"c0",x"79"),
  1757 => (x"49",x"66",x"c4",x"c1"),
  1758 => (x"c1",x"81",x"d4",x"c1"),
  1759 => (x"c1",x"4a",x"66",x"c4"),
  1760 => (x"ca",x"c1",x"82",x"d8"),
  1761 => (x"d8",x"c1",x"7a",x"f4"),
  1762 => (x"c4",x"c1",x"79",x"fc"),
  1763 => (x"e0",x"c1",x"49",x"66"),
  1764 => (x"e3",x"dc",x"c1",x"81"),
  1765 => (x"d8",x"d0",x"ff",x"79"),
  1766 => (x"48",x"66",x"d0",x"87"),
  1767 => (x"26",x"8e",x"cc",x"ff"),
  1768 => (x"26",x"4c",x"26",x"4d"),
  1769 => (x"1e",x"4f",x"26",x"4b"),
  1770 => (x"f5",x"c2",x"1e",x"c7"),
  1771 => (x"c1",x"1e",x"bf",x"d8"),
  1772 => (x"c2",x"1e",x"e0",x"f1"),
  1773 => (x"bf",x"97",x"c8",x"f4"),
  1774 => (x"87",x"f9",x"ee",x"49"),
  1775 => (x"49",x"e0",x"f1",x"c1"),
  1776 => (x"87",x"f6",x"e0",x"c0"),
  1777 => (x"4f",x"26",x"8e",x"f4"),
  1778 => (x"d4",x"f1",x"c1",x"1e"),
  1779 => (x"c1",x"50",x"c0",x"48"),
  1780 => (x"49",x"bf",x"cc",x"f3"),
  1781 => (x"87",x"ce",x"d5",x"ff"),
  1782 => (x"4f",x"26",x"48",x"c0"),
  1783 => (x"c7",x"1e",x"73",x"1e"),
  1784 => (x"f5",x"c2",x"87",x"cc"),
  1785 => (x"50",x"c0",x"48",x"e4"),
  1786 => (x"c3",x"48",x"d4",x"ff"),
  1787 => (x"ca",x"c1",x"78",x"ff"),
  1788 => (x"d7",x"fe",x"49",x"fc"),
  1789 => (x"e2",x"fe",x"87",x"d3"),
  1790 => (x"98",x"70",x"87",x"e6"),
  1791 => (x"fe",x"87",x"cd",x"02"),
  1792 => (x"70",x"87",x"c4",x"ec"),
  1793 => (x"87",x"c4",x"02",x"98"),
  1794 => (x"87",x"c2",x"4a",x"c1"),
  1795 => (x"9a",x"72",x"4a",x"c0"),
  1796 => (x"c1",x"87",x"c8",x"02"),
  1797 => (x"fe",x"49",x"c8",x"cb"),
  1798 => (x"c2",x"87",x"ee",x"d6"),
  1799 => (x"c0",x"48",x"d8",x"f5"),
  1800 => (x"c8",x"f4",x"c2",x"78"),
  1801 => (x"49",x"50",x"c0",x"48"),
  1802 => (x"fe",x"87",x"fc",x"fd"),
  1803 => (x"4b",x"70",x"87",x"da"),
  1804 => (x"87",x"ce",x"02",x"9b"),
  1805 => (x"5b",x"fc",x"f2",x"c1"),
  1806 => (x"ef",x"dd",x"49",x"c7"),
  1807 => (x"df",x"49",x"c1",x"87"),
  1808 => (x"f2",x"c2",x"87",x"cb"),
  1809 => (x"d1",x"e0",x"c0",x"87"),
  1810 => (x"e3",x"ee",x"c0",x"87"),
  1811 => (x"87",x"f5",x"ff",x"87"),
  1812 => (x"4f",x"26",x"4b",x"26"),
  1813 => (x"00",x"00",x"00",x"00"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"00",x"00",x"00",x"01"),
  1816 => (x"00",x"00",x"13",x"1e"),
  1817 => (x"00",x"00",x"2d",x"70"),
  1818 => (x"54",x"00",x"00",x"00"),
  1819 => (x"00",x"00",x"13",x"1e"),
  1820 => (x"00",x"00",x"2d",x"8e"),
  1821 => (x"54",x"00",x"00",x"00"),
  1822 => (x"00",x"00",x"13",x"1e"),
  1823 => (x"00",x"00",x"2d",x"ac"),
  1824 => (x"54",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"13",x"1e"),
  1826 => (x"00",x"00",x"2d",x"ca"),
  1827 => (x"54",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"13",x"1e"),
  1829 => (x"00",x"00",x"2d",x"e8"),
  1830 => (x"54",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"13",x"1e"),
  1832 => (x"00",x"00",x"2e",x"06"),
  1833 => (x"54",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"13",x"1e"),
  1835 => (x"00",x"00",x"2e",x"24"),
  1836 => (x"54",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"16",x"45"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"54",x"00",x"00",x"00"),
  1840 => (x"00",x"00",x"13",x"f7"),
  1841 => (x"00",x"00",x"00",x"00"),
  1842 => (x"54",x"00",x"00",x"00"),
  1843 => (x"00",x"00",x"12",x"cc"),
  1844 => (x"db",x"86",x"fc",x"1e"),
  1845 => (x"fc",x"7e",x"70",x"87"),
  1846 => (x"1e",x"4f",x"26",x"8e"),
  1847 => (x"c0",x"48",x"f0",x"fe"),
  1848 => (x"79",x"09",x"cd",x"78"),
  1849 => (x"1e",x"4f",x"26",x"09"),
  1850 => (x"49",x"d0",x"f3",x"c1"),
  1851 => (x"4f",x"26",x"87",x"ed"),
  1852 => (x"bf",x"f0",x"fe",x"1e"),
  1853 => (x"1e",x"4f",x"26",x"48"),
  1854 => (x"c1",x"48",x"f0",x"fe"),
  1855 => (x"1e",x"4f",x"26",x"78"),
  1856 => (x"c0",x"48",x"f0",x"fe"),
  1857 => (x"1e",x"4f",x"26",x"78"),
  1858 => (x"52",x"c0",x"4a",x"71"),
  1859 => (x"0e",x"4f",x"26",x"51"),
  1860 => (x"5d",x"5c",x"5b",x"5e"),
  1861 => (x"71",x"86",x"f4",x"0e"),
  1862 => (x"7e",x"6d",x"97",x"4d"),
  1863 => (x"97",x"4c",x"a5",x"c1"),
  1864 => (x"a6",x"c8",x"48",x"6c"),
  1865 => (x"c4",x"48",x"6e",x"58"),
  1866 => (x"c5",x"05",x"a8",x"66"),
  1867 => (x"c0",x"48",x"ff",x"87"),
  1868 => (x"ca",x"ff",x"87",x"e6"),
  1869 => (x"49",x"a5",x"c2",x"87"),
  1870 => (x"71",x"4b",x"6c",x"97"),
  1871 => (x"6b",x"97",x"4b",x"a3"),
  1872 => (x"7e",x"6c",x"97",x"4b"),
  1873 => (x"80",x"c1",x"48",x"6e"),
  1874 => (x"c7",x"58",x"a6",x"c8"),
  1875 => (x"58",x"a6",x"cc",x"98"),
  1876 => (x"fe",x"7c",x"97",x"70"),
  1877 => (x"48",x"73",x"87",x"e1"),
  1878 => (x"4d",x"26",x"8e",x"f4"),
  1879 => (x"4b",x"26",x"4c",x"26"),
  1880 => (x"73",x"1e",x"4f",x"26"),
  1881 => (x"fe",x"86",x"f4",x"1e"),
  1882 => (x"bf",x"e0",x"87",x"d5"),
  1883 => (x"e0",x"c0",x"49",x"4b"),
  1884 => (x"c0",x"02",x"99",x"c0"),
  1885 => (x"4a",x"73",x"87",x"ea"),
  1886 => (x"c2",x"9a",x"ff",x"c3"),
  1887 => (x"bf",x"97",x"d8",x"f9"),
  1888 => (x"da",x"f9",x"c2",x"49"),
  1889 => (x"c2",x"51",x"72",x"81"),
  1890 => (x"bf",x"97",x"d8",x"f9"),
  1891 => (x"c1",x"48",x"6e",x"7e"),
  1892 => (x"58",x"a6",x"c8",x"80"),
  1893 => (x"a6",x"cc",x"98",x"c7"),
  1894 => (x"d8",x"f9",x"c2",x"58"),
  1895 => (x"50",x"66",x"c8",x"48"),
  1896 => (x"70",x"87",x"cd",x"fd"),
  1897 => (x"87",x"cf",x"fd",x"7e"),
  1898 => (x"4b",x"26",x"8e",x"f4"),
  1899 => (x"c2",x"1e",x"4f",x"26"),
  1900 => (x"fd",x"49",x"d8",x"f9"),
  1901 => (x"f5",x"c1",x"87",x"d1"),
  1902 => (x"de",x"fc",x"49",x"e2"),
  1903 => (x"87",x"f0",x"c3",x"87"),
  1904 => (x"73",x"1e",x"4f",x"26"),
  1905 => (x"d8",x"f9",x"c2",x"1e"),
  1906 => (x"87",x"c3",x"fd",x"49"),
  1907 => (x"b7",x"c0",x"4a",x"70"),
  1908 => (x"cc",x"c2",x"04",x"aa"),
  1909 => (x"aa",x"f0",x"c3",x"87"),
  1910 => (x"c1",x"87",x"c9",x"05"),
  1911 => (x"c1",x"48",x"e8",x"f9"),
  1912 => (x"87",x"ed",x"c1",x"78"),
  1913 => (x"05",x"aa",x"e0",x"c3"),
  1914 => (x"f9",x"c1",x"87",x"c9"),
  1915 => (x"78",x"c1",x"48",x"ec"),
  1916 => (x"c1",x"87",x"de",x"c1"),
  1917 => (x"02",x"bf",x"ec",x"f9"),
  1918 => (x"c0",x"c2",x"87",x"c6"),
  1919 => (x"87",x"c2",x"4b",x"a2"),
  1920 => (x"f9",x"c1",x"4b",x"72"),
  1921 => (x"c0",x"02",x"bf",x"e8"),
  1922 => (x"49",x"73",x"87",x"e0"),
  1923 => (x"91",x"29",x"b7",x"c4"),
  1924 => (x"81",x"f0",x"f9",x"c1"),
  1925 => (x"9a",x"cf",x"4a",x"73"),
  1926 => (x"48",x"c1",x"92",x"c2"),
  1927 => (x"4a",x"70",x"30",x"72"),
  1928 => (x"48",x"72",x"ba",x"ff"),
  1929 => (x"79",x"70",x"98",x"69"),
  1930 => (x"49",x"73",x"87",x"db"),
  1931 => (x"91",x"29",x"b7",x"c4"),
  1932 => (x"81",x"f0",x"f9",x"c1"),
  1933 => (x"9a",x"cf",x"4a",x"73"),
  1934 => (x"48",x"c3",x"92",x"c2"),
  1935 => (x"4a",x"70",x"30",x"72"),
  1936 => (x"70",x"b0",x"69",x"48"),
  1937 => (x"ec",x"f9",x"c1",x"79"),
  1938 => (x"c1",x"78",x"c0",x"48"),
  1939 => (x"c0",x"48",x"e8",x"f9"),
  1940 => (x"d8",x"f9",x"c2",x"78"),
  1941 => (x"87",x"f7",x"fa",x"49"),
  1942 => (x"b7",x"c0",x"4a",x"70"),
  1943 => (x"f4",x"fd",x"03",x"aa"),
  1944 => (x"26",x"48",x"c0",x"87"),
  1945 => (x"00",x"4f",x"26",x"4b"),
  1946 => (x"00",x"00",x"00",x"00"),
  1947 => (x"00",x"00",x"00",x"00"),
  1948 => (x"00",x"00",x"00",x"00"),
  1949 => (x"84",x"84",x"84",x"84"),
  1950 => (x"84",x"84",x"84",x"84"),
  1951 => (x"84",x"84",x"84",x"84"),
  1952 => (x"84",x"84",x"84",x"84"),
  1953 => (x"84",x"84",x"84",x"84"),
  1954 => (x"84",x"84",x"84",x"84"),
  1955 => (x"84",x"84",x"84",x"84"),
  1956 => (x"84",x"84",x"84",x"84"),
  1957 => (x"84",x"84",x"84",x"84"),
  1958 => (x"84",x"84",x"84",x"84"),
  1959 => (x"84",x"84",x"84",x"84"),
  1960 => (x"84",x"84",x"84",x"84"),
  1961 => (x"84",x"84",x"84",x"84"),
  1962 => (x"84",x"84",x"84",x"84"),
  1963 => (x"84",x"84",x"84",x"84"),
  1964 => (x"72",x"4a",x"c0",x"1e"),
  1965 => (x"c1",x"91",x"c4",x"49"),
  1966 => (x"c0",x"81",x"f0",x"f9"),
  1967 => (x"d0",x"82",x"c1",x"79"),
  1968 => (x"ee",x"04",x"aa",x"b7"),
  1969 => (x"0e",x"4f",x"26",x"87"),
  1970 => (x"5d",x"5c",x"5b",x"5e"),
  1971 => (x"f8",x"4d",x"71",x"0e"),
  1972 => (x"4a",x"75",x"87",x"ed"),
  1973 => (x"92",x"2a",x"b7",x"c4"),
  1974 => (x"82",x"f0",x"f9",x"c1"),
  1975 => (x"9c",x"cf",x"4c",x"75"),
  1976 => (x"49",x"6a",x"94",x"c2"),
  1977 => (x"c3",x"2b",x"74",x"4b"),
  1978 => (x"74",x"48",x"c2",x"9b"),
  1979 => (x"ff",x"4c",x"70",x"30"),
  1980 => (x"71",x"48",x"74",x"bc"),
  1981 => (x"f7",x"7a",x"70",x"98"),
  1982 => (x"48",x"73",x"87",x"fd"),
  1983 => (x"4c",x"26",x"4d",x"26"),
  1984 => (x"4f",x"26",x"4b",x"26"),
  1985 => (x"48",x"d0",x"ff",x"1e"),
  1986 => (x"71",x"78",x"e1",x"c8"),
  1987 => (x"08",x"d4",x"ff",x"48"),
  1988 => (x"1e",x"4f",x"26",x"78"),
  1989 => (x"c8",x"48",x"d0",x"ff"),
  1990 => (x"48",x"71",x"78",x"e1"),
  1991 => (x"78",x"08",x"d4",x"ff"),
  1992 => (x"ff",x"48",x"66",x"c4"),
  1993 => (x"26",x"78",x"08",x"d4"),
  1994 => (x"4a",x"71",x"1e",x"4f"),
  1995 => (x"1e",x"49",x"66",x"c4"),
  1996 => (x"de",x"ff",x"49",x"72"),
  1997 => (x"48",x"d0",x"ff",x"87"),
  1998 => (x"fc",x"78",x"e0",x"c0"),
  1999 => (x"1e",x"4f",x"26",x"8e"),
  2000 => (x"4b",x"71",x"1e",x"73"),
  2001 => (x"1e",x"49",x"66",x"c8"),
  2002 => (x"e0",x"c1",x"4a",x"73"),
  2003 => (x"d8",x"ff",x"49",x"a2"),
  2004 => (x"26",x"8e",x"fc",x"87"),
  2005 => (x"1e",x"4f",x"26",x"4b"),
  2006 => (x"c8",x"48",x"d0",x"ff"),
  2007 => (x"48",x"71",x"78",x"c9"),
  2008 => (x"78",x"08",x"d4",x"ff"),
  2009 => (x"71",x"1e",x"4f",x"26"),
  2010 => (x"87",x"eb",x"49",x"4a"),
  2011 => (x"c8",x"48",x"d0",x"ff"),
  2012 => (x"1e",x"4f",x"26",x"78"),
  2013 => (x"4b",x"71",x"1e",x"73"),
  2014 => (x"bf",x"f0",x"f9",x"c2"),
  2015 => (x"c2",x"87",x"c3",x"02"),
  2016 => (x"d0",x"ff",x"87",x"eb"),
  2017 => (x"78",x"c9",x"c8",x"48"),
  2018 => (x"e0",x"c0",x"48",x"73"),
  2019 => (x"08",x"d4",x"ff",x"b0"),
  2020 => (x"e4",x"f9",x"c2",x"78"),
  2021 => (x"c8",x"78",x"c0",x"48"),
  2022 => (x"87",x"c5",x"02",x"66"),
  2023 => (x"c2",x"49",x"ff",x"c3"),
  2024 => (x"c2",x"49",x"c0",x"87"),
  2025 => (x"cc",x"59",x"ec",x"f9"),
  2026 => (x"87",x"c6",x"02",x"66"),
  2027 => (x"4a",x"d5",x"d5",x"c5"),
  2028 => (x"ff",x"cf",x"87",x"c4"),
  2029 => (x"f9",x"c2",x"4a",x"ff"),
  2030 => (x"f9",x"c2",x"5a",x"f0"),
  2031 => (x"78",x"c1",x"48",x"f0"),
  2032 => (x"4f",x"26",x"4b",x"26"),
  2033 => (x"5c",x"5b",x"5e",x"0e"),
  2034 => (x"4d",x"71",x"0e",x"5d"),
  2035 => (x"bf",x"ec",x"f9",x"c2"),
  2036 => (x"02",x"9d",x"75",x"4b"),
  2037 => (x"c8",x"49",x"87",x"cb"),
  2038 => (x"ec",x"fd",x"c1",x"91"),
  2039 => (x"c4",x"82",x"71",x"4a"),
  2040 => (x"ec",x"c1",x"c2",x"87"),
  2041 => (x"12",x"4c",x"c0",x"4a"),
  2042 => (x"c2",x"99",x"73",x"49"),
  2043 => (x"48",x"bf",x"e8",x"f9"),
  2044 => (x"d4",x"ff",x"b8",x"71"),
  2045 => (x"b7",x"c1",x"78",x"08"),
  2046 => (x"b7",x"c8",x"84",x"2b"),
  2047 => (x"87",x"e7",x"04",x"ac"),
  2048 => (x"bf",x"e4",x"f9",x"c2"),
  2049 => (x"c2",x"80",x"c8",x"48"),
  2050 => (x"26",x"58",x"e8",x"f9"),
  2051 => (x"26",x"4c",x"26",x"4d"),
  2052 => (x"1e",x"4f",x"26",x"4b"),
  2053 => (x"4b",x"71",x"1e",x"73"),
  2054 => (x"02",x"9a",x"4a",x"13"),
  2055 => (x"49",x"72",x"87",x"cb"),
  2056 => (x"13",x"87",x"e1",x"fe"),
  2057 => (x"f5",x"05",x"9a",x"4a"),
  2058 => (x"26",x"4b",x"26",x"87"),
  2059 => (x"f9",x"c2",x"1e",x"4f"),
  2060 => (x"c2",x"49",x"bf",x"e4"),
  2061 => (x"c1",x"48",x"e4",x"f9"),
  2062 => (x"c0",x"c4",x"78",x"a1"),
  2063 => (x"db",x"03",x"a9",x"b7"),
  2064 => (x"48",x"d4",x"ff",x"87"),
  2065 => (x"bf",x"e8",x"f9",x"c2"),
  2066 => (x"e4",x"f9",x"c2",x"78"),
  2067 => (x"f9",x"c2",x"49",x"bf"),
  2068 => (x"a1",x"c1",x"48",x"e4"),
  2069 => (x"b7",x"c0",x"c4",x"78"),
  2070 => (x"87",x"e5",x"04",x"a9"),
  2071 => (x"c8",x"48",x"d0",x"ff"),
  2072 => (x"f0",x"f9",x"c2",x"78"),
  2073 => (x"26",x"78",x"c0",x"48"),
  2074 => (x"00",x"00",x"00",x"4f"),
  2075 => (x"00",x"00",x"00",x"00"),
  2076 => (x"00",x"00",x"00",x"00"),
  2077 => (x"5f",x"00",x"00",x"00"),
  2078 => (x"00",x"00",x"00",x"5f"),
  2079 => (x"00",x"03",x"03",x"00"),
  2080 => (x"00",x"00",x"03",x"03"),
  2081 => (x"14",x"7f",x"7f",x"14"),
  2082 => (x"00",x"14",x"7f",x"7f"),
  2083 => (x"6b",x"2e",x"24",x"00"),
  2084 => (x"00",x"12",x"3a",x"6b"),
  2085 => (x"18",x"36",x"6a",x"4c"),
  2086 => (x"00",x"32",x"56",x"6c"),
  2087 => (x"59",x"4f",x"7e",x"30"),
  2088 => (x"40",x"68",x"3a",x"77"),
  2089 => (x"07",x"04",x"00",x"00"),
  2090 => (x"00",x"00",x"00",x"03"),
  2091 => (x"3e",x"1c",x"00",x"00"),
  2092 => (x"00",x"00",x"41",x"63"),
  2093 => (x"63",x"41",x"00",x"00"),
  2094 => (x"00",x"00",x"1c",x"3e"),
  2095 => (x"1c",x"3e",x"2a",x"08"),
  2096 => (x"08",x"2a",x"3e",x"1c"),
  2097 => (x"3e",x"08",x"08",x"00"),
  2098 => (x"00",x"08",x"08",x"3e"),
  2099 => (x"e0",x"80",x"00",x"00"),
  2100 => (x"00",x"00",x"00",x"60"),
  2101 => (x"08",x"08",x"08",x"00"),
  2102 => (x"00",x"08",x"08",x"08"),
  2103 => (x"60",x"00",x"00",x"00"),
  2104 => (x"00",x"00",x"00",x"60"),
  2105 => (x"18",x"30",x"60",x"40"),
  2106 => (x"01",x"03",x"06",x"0c"),
  2107 => (x"59",x"7f",x"3e",x"00"),
  2108 => (x"00",x"3e",x"7f",x"4d"),
  2109 => (x"7f",x"06",x"04",x"00"),
  2110 => (x"00",x"00",x"00",x"7f"),
  2111 => (x"71",x"63",x"42",x"00"),
  2112 => (x"00",x"46",x"4f",x"59"),
  2113 => (x"49",x"63",x"22",x"00"),
  2114 => (x"00",x"36",x"7f",x"49"),
  2115 => (x"13",x"16",x"1c",x"18"),
  2116 => (x"00",x"10",x"7f",x"7f"),
  2117 => (x"45",x"67",x"27",x"00"),
  2118 => (x"00",x"39",x"7d",x"45"),
  2119 => (x"4b",x"7e",x"3c",x"00"),
  2120 => (x"00",x"30",x"79",x"49"),
  2121 => (x"71",x"01",x"01",x"00"),
  2122 => (x"00",x"07",x"0f",x"79"),
  2123 => (x"49",x"7f",x"36",x"00"),
  2124 => (x"00",x"36",x"7f",x"49"),
  2125 => (x"49",x"4f",x"06",x"00"),
  2126 => (x"00",x"1e",x"3f",x"69"),
  2127 => (x"66",x"00",x"00",x"00"),
  2128 => (x"00",x"00",x"00",x"66"),
  2129 => (x"e6",x"80",x"00",x"00"),
  2130 => (x"00",x"00",x"00",x"66"),
  2131 => (x"14",x"08",x"08",x"00"),
  2132 => (x"00",x"22",x"22",x"14"),
  2133 => (x"14",x"14",x"14",x"00"),
  2134 => (x"00",x"14",x"14",x"14"),
  2135 => (x"14",x"22",x"22",x"00"),
  2136 => (x"00",x"08",x"08",x"14"),
  2137 => (x"51",x"03",x"02",x"00"),
  2138 => (x"00",x"06",x"0f",x"59"),
  2139 => (x"5d",x"41",x"7f",x"3e"),
  2140 => (x"00",x"1e",x"1f",x"55"),
  2141 => (x"09",x"7f",x"7e",x"00"),
  2142 => (x"00",x"7e",x"7f",x"09"),
  2143 => (x"49",x"7f",x"7f",x"00"),
  2144 => (x"00",x"36",x"7f",x"49"),
  2145 => (x"63",x"3e",x"1c",x"00"),
  2146 => (x"00",x"41",x"41",x"41"),
  2147 => (x"41",x"7f",x"7f",x"00"),
  2148 => (x"00",x"1c",x"3e",x"63"),
  2149 => (x"49",x"7f",x"7f",x"00"),
  2150 => (x"00",x"41",x"41",x"49"),
  2151 => (x"09",x"7f",x"7f",x"00"),
  2152 => (x"00",x"01",x"01",x"09"),
  2153 => (x"41",x"7f",x"3e",x"00"),
  2154 => (x"00",x"7a",x"7b",x"49"),
  2155 => (x"08",x"7f",x"7f",x"00"),
  2156 => (x"00",x"7f",x"7f",x"08"),
  2157 => (x"7f",x"41",x"00",x"00"),
  2158 => (x"00",x"00",x"41",x"7f"),
  2159 => (x"40",x"60",x"20",x"00"),
  2160 => (x"00",x"3f",x"7f",x"40"),
  2161 => (x"1c",x"08",x"7f",x"7f"),
  2162 => (x"00",x"41",x"63",x"36"),
  2163 => (x"40",x"7f",x"7f",x"00"),
  2164 => (x"00",x"40",x"40",x"40"),
  2165 => (x"0c",x"06",x"7f",x"7f"),
  2166 => (x"00",x"7f",x"7f",x"06"),
  2167 => (x"0c",x"06",x"7f",x"7f"),
  2168 => (x"00",x"7f",x"7f",x"18"),
  2169 => (x"41",x"7f",x"3e",x"00"),
  2170 => (x"00",x"3e",x"7f",x"41"),
  2171 => (x"09",x"7f",x"7f",x"00"),
  2172 => (x"00",x"06",x"0f",x"09"),
  2173 => (x"61",x"41",x"7f",x"3e"),
  2174 => (x"00",x"40",x"7e",x"7f"),
  2175 => (x"09",x"7f",x"7f",x"00"),
  2176 => (x"00",x"66",x"7f",x"19"),
  2177 => (x"4d",x"6f",x"26",x"00"),
  2178 => (x"00",x"32",x"7b",x"59"),
  2179 => (x"7f",x"01",x"01",x"00"),
  2180 => (x"00",x"01",x"01",x"7f"),
  2181 => (x"40",x"7f",x"3f",x"00"),
  2182 => (x"00",x"3f",x"7f",x"40"),
  2183 => (x"70",x"3f",x"0f",x"00"),
  2184 => (x"00",x"0f",x"3f",x"70"),
  2185 => (x"18",x"30",x"7f",x"7f"),
  2186 => (x"00",x"7f",x"7f",x"30"),
  2187 => (x"1c",x"36",x"63",x"41"),
  2188 => (x"41",x"63",x"36",x"1c"),
  2189 => (x"7c",x"06",x"03",x"01"),
  2190 => (x"01",x"03",x"06",x"7c"),
  2191 => (x"4d",x"59",x"71",x"61"),
  2192 => (x"00",x"41",x"43",x"47"),
  2193 => (x"7f",x"7f",x"00",x"00"),
  2194 => (x"00",x"00",x"41",x"41"),
  2195 => (x"0c",x"06",x"03",x"01"),
  2196 => (x"40",x"60",x"30",x"18"),
  2197 => (x"41",x"41",x"00",x"00"),
  2198 => (x"00",x"00",x"7f",x"7f"),
  2199 => (x"03",x"06",x"0c",x"08"),
  2200 => (x"00",x"08",x"0c",x"06"),
  2201 => (x"80",x"80",x"80",x"80"),
  2202 => (x"00",x"80",x"80",x"80"),
  2203 => (x"03",x"00",x"00",x"00"),
  2204 => (x"00",x"00",x"04",x"07"),
  2205 => (x"54",x"74",x"20",x"00"),
  2206 => (x"00",x"78",x"7c",x"54"),
  2207 => (x"44",x"7f",x"7f",x"00"),
  2208 => (x"00",x"38",x"7c",x"44"),
  2209 => (x"44",x"7c",x"38",x"00"),
  2210 => (x"00",x"00",x"44",x"44"),
  2211 => (x"44",x"7c",x"38",x"00"),
  2212 => (x"00",x"7f",x"7f",x"44"),
  2213 => (x"54",x"7c",x"38",x"00"),
  2214 => (x"00",x"18",x"5c",x"54"),
  2215 => (x"7f",x"7e",x"04",x"00"),
  2216 => (x"00",x"00",x"05",x"05"),
  2217 => (x"a4",x"bc",x"18",x"00"),
  2218 => (x"00",x"7c",x"fc",x"a4"),
  2219 => (x"04",x"7f",x"7f",x"00"),
  2220 => (x"00",x"78",x"7c",x"04"),
  2221 => (x"3d",x"00",x"00",x"00"),
  2222 => (x"00",x"00",x"40",x"7d"),
  2223 => (x"80",x"80",x"80",x"00"),
  2224 => (x"00",x"00",x"7d",x"fd"),
  2225 => (x"10",x"7f",x"7f",x"00"),
  2226 => (x"00",x"44",x"6c",x"38"),
  2227 => (x"3f",x"00",x"00",x"00"),
  2228 => (x"00",x"00",x"40",x"7f"),
  2229 => (x"18",x"0c",x"7c",x"7c"),
  2230 => (x"00",x"78",x"7c",x"0c"),
  2231 => (x"04",x"7c",x"7c",x"00"),
  2232 => (x"00",x"78",x"7c",x"04"),
  2233 => (x"44",x"7c",x"38",x"00"),
  2234 => (x"00",x"38",x"7c",x"44"),
  2235 => (x"24",x"fc",x"fc",x"00"),
  2236 => (x"00",x"18",x"3c",x"24"),
  2237 => (x"24",x"3c",x"18",x"00"),
  2238 => (x"00",x"fc",x"fc",x"24"),
  2239 => (x"04",x"7c",x"7c",x"00"),
  2240 => (x"00",x"08",x"0c",x"04"),
  2241 => (x"54",x"5c",x"48",x"00"),
  2242 => (x"00",x"20",x"74",x"54"),
  2243 => (x"7f",x"3f",x"04",x"00"),
  2244 => (x"00",x"00",x"44",x"44"),
  2245 => (x"40",x"7c",x"3c",x"00"),
  2246 => (x"00",x"7c",x"7c",x"40"),
  2247 => (x"60",x"3c",x"1c",x"00"),
  2248 => (x"00",x"1c",x"3c",x"60"),
  2249 => (x"30",x"60",x"7c",x"3c"),
  2250 => (x"00",x"3c",x"7c",x"60"),
  2251 => (x"10",x"38",x"6c",x"44"),
  2252 => (x"00",x"44",x"6c",x"38"),
  2253 => (x"e0",x"bc",x"1c",x"00"),
  2254 => (x"00",x"1c",x"3c",x"60"),
  2255 => (x"74",x"64",x"44",x"00"),
  2256 => (x"00",x"44",x"4c",x"5c"),
  2257 => (x"3e",x"08",x"08",x"00"),
  2258 => (x"00",x"41",x"41",x"77"),
  2259 => (x"7f",x"00",x"00",x"00"),
  2260 => (x"00",x"00",x"00",x"7f"),
  2261 => (x"77",x"41",x"41",x"00"),
  2262 => (x"00",x"08",x"08",x"3e"),
  2263 => (x"03",x"01",x"01",x"02"),
  2264 => (x"00",x"01",x"02",x"02"),
  2265 => (x"7f",x"7f",x"7f",x"7f"),
  2266 => (x"00",x"7f",x"7f",x"7f"),
  2267 => (x"1c",x"1c",x"08",x"08"),
  2268 => (x"7f",x"7f",x"3e",x"3e"),
  2269 => (x"3e",x"3e",x"7f",x"7f"),
  2270 => (x"08",x"08",x"1c",x"1c"),
  2271 => (x"7c",x"18",x"10",x"00"),
  2272 => (x"00",x"10",x"18",x"7c"),
  2273 => (x"7c",x"30",x"10",x"00"),
  2274 => (x"00",x"10",x"30",x"7c"),
  2275 => (x"60",x"60",x"30",x"10"),
  2276 => (x"00",x"06",x"1e",x"78"),
  2277 => (x"18",x"3c",x"66",x"42"),
  2278 => (x"00",x"42",x"66",x"3c"),
  2279 => (x"c2",x"6a",x"38",x"78"),
  2280 => (x"00",x"38",x"6c",x"c6"),
  2281 => (x"60",x"00",x"00",x"60"),
  2282 => (x"00",x"60",x"00",x"00"),
  2283 => (x"5c",x"5b",x"5e",x"0e"),
  2284 => (x"86",x"fc",x"0e",x"5d"),
  2285 => (x"f9",x"c2",x"7e",x"71"),
  2286 => (x"c0",x"4c",x"bf",x"f8"),
  2287 => (x"c4",x"1e",x"c0",x"4b"),
  2288 => (x"c4",x"02",x"ab",x"66"),
  2289 => (x"c2",x"4d",x"c0",x"87"),
  2290 => (x"75",x"4d",x"c1",x"87"),
  2291 => (x"ee",x"49",x"73",x"1e"),
  2292 => (x"86",x"c8",x"87",x"e1"),
  2293 => (x"ef",x"49",x"e0",x"c0"),
  2294 => (x"a4",x"c4",x"87",x"ea"),
  2295 => (x"f0",x"49",x"6a",x"4a"),
  2296 => (x"c8",x"f1",x"87",x"f1"),
  2297 => (x"c1",x"84",x"cc",x"87"),
  2298 => (x"ab",x"b7",x"c8",x"83"),
  2299 => (x"87",x"cd",x"ff",x"04"),
  2300 => (x"4d",x"26",x"8e",x"fc"),
  2301 => (x"4b",x"26",x"4c",x"26"),
  2302 => (x"71",x"1e",x"4f",x"26"),
  2303 => (x"fc",x"f9",x"c2",x"4a"),
  2304 => (x"fc",x"f9",x"c2",x"5a"),
  2305 => (x"49",x"78",x"c7",x"48"),
  2306 => (x"26",x"87",x"e1",x"fe"),
  2307 => (x"1e",x"73",x"1e",x"4f"),
  2308 => (x"0b",x"fc",x"4b",x"71"),
  2309 => (x"4a",x"73",x"0b",x"7b"),
  2310 => (x"c0",x"c1",x"9a",x"c1"),
  2311 => (x"c5",x"ed",x"49",x"a2"),
  2312 => (x"fc",x"dd",x"c2",x"87"),
  2313 => (x"26",x"4b",x"26",x"5b"),
  2314 => (x"4a",x"71",x"1e",x"4f"),
  2315 => (x"72",x"1e",x"66",x"c4"),
  2316 => (x"87",x"cb",x"ec",x"49"),
  2317 => (x"4f",x"26",x"8e",x"fc"),
  2318 => (x"48",x"d4",x"ff",x"1e"),
  2319 => (x"ff",x"78",x"ff",x"c3"),
  2320 => (x"e1",x"c0",x"48",x"d0"),
  2321 => (x"48",x"d4",x"ff",x"78"),
  2322 => (x"48",x"71",x"78",x"c1"),
  2323 => (x"d4",x"ff",x"30",x"c4"),
  2324 => (x"d0",x"ff",x"78",x"08"),
  2325 => (x"78",x"e0",x"c0",x"48"),
  2326 => (x"5e",x"0e",x"4f",x"26"),
  2327 => (x"0e",x"5d",x"5c",x"5b"),
  2328 => (x"a6",x"c8",x"86",x"ec"),
  2329 => (x"c4",x"78",x"c0",x"48"),
  2330 => (x"78",x"bf",x"ec",x"80"),
  2331 => (x"f9",x"c2",x"80",x"f8"),
  2332 => (x"c2",x"78",x"bf",x"f8"),
  2333 => (x"4c",x"bf",x"c0",x"fa"),
  2334 => (x"c2",x"4d",x"bf",x"e8"),
  2335 => (x"49",x"bf",x"f8",x"dd"),
  2336 => (x"c7",x"87",x"ff",x"e4"),
  2337 => (x"87",x"ff",x"e8",x"49"),
  2338 => (x"99",x"c2",x"49",x"70"),
  2339 => (x"c2",x"87",x"d0",x"05"),
  2340 => (x"49",x"bf",x"f0",x"dd"),
  2341 => (x"66",x"cc",x"b9",x"ff"),
  2342 => (x"02",x"99",x"c1",x"99"),
  2343 => (x"c8",x"87",x"cb",x"c2"),
  2344 => (x"c8",x"ff",x"48",x"a6"),
  2345 => (x"49",x"c7",x"78",x"bf"),
  2346 => (x"70",x"87",x"dc",x"e8"),
  2347 => (x"71",x"7e",x"74",x"49"),
  2348 => (x"87",x"cd",x"05",x"99"),
  2349 => (x"c1",x"49",x"66",x"cc"),
  2350 => (x"71",x"7e",x"74",x"99"),
  2351 => (x"c4",x"c1",x"02",x"99"),
  2352 => (x"4c",x"c8",x"ff",x"87"),
  2353 => (x"cc",x"4b",x"66",x"c8"),
  2354 => (x"bf",x"ec",x"48",x"a6"),
  2355 => (x"87",x"f2",x"e3",x"78"),
  2356 => (x"6c",x"5b",x"a6",x"cc"),
  2357 => (x"d4",x"88",x"73",x"48"),
  2358 => (x"e8",x"cf",x"58",x"a6"),
  2359 => (x"87",x"d1",x"06",x"a8"),
  2360 => (x"bf",x"ec",x"dd",x"c2"),
  2361 => (x"c2",x"b9",x"c1",x"49"),
  2362 => (x"71",x"59",x"f0",x"dd"),
  2363 => (x"6c",x"87",x"c9",x"fd"),
  2364 => (x"e7",x"49",x"c7",x"4b"),
  2365 => (x"98",x"70",x"87",x"d1"),
  2366 => (x"87",x"cb",x"ff",x"05"),
  2367 => (x"c1",x"49",x"66",x"cc"),
  2368 => (x"c2",x"ff",x"05",x"99"),
  2369 => (x"c2",x"4c",x"6e",x"87"),
  2370 => (x"4a",x"bf",x"f8",x"dd"),
  2371 => (x"dd",x"c2",x"ba",x"c1"),
  2372 => (x"0a",x"fc",x"5a",x"fc"),
  2373 => (x"9a",x"c1",x"0a",x"7a"),
  2374 => (x"49",x"a2",x"c0",x"c1"),
  2375 => (x"c1",x"87",x"c7",x"e9"),
  2376 => (x"e2",x"e6",x"49",x"da"),
  2377 => (x"48",x"a6",x"c8",x"87"),
  2378 => (x"dd",x"c2",x"78",x"c1"),
  2379 => (x"66",x"cc",x"48",x"f0"),
  2380 => (x"f8",x"dd",x"c2",x"78"),
  2381 => (x"c7",x"c1",x"05",x"bf"),
  2382 => (x"c0",x"c0",x"c8",x"87"),
  2383 => (x"dc",x"dd",x"c2",x"4b"),
  2384 => (x"14",x"4c",x"6e",x"7e"),
  2385 => (x"87",x"ff",x"e5",x"49"),
  2386 => (x"c0",x"02",x"98",x"70"),
  2387 => (x"b5",x"73",x"87",x"c2"),
  2388 => (x"05",x"2b",x"b7",x"c1"),
  2389 => (x"75",x"87",x"ec",x"ff"),
  2390 => (x"99",x"ff",x"c3",x"49"),
  2391 => (x"49",x"c0",x"1e",x"71"),
  2392 => (x"75",x"87",x"c6",x"fb"),
  2393 => (x"29",x"b7",x"c8",x"49"),
  2394 => (x"49",x"c1",x"1e",x"71"),
  2395 => (x"c8",x"87",x"fa",x"fa"),
  2396 => (x"49",x"fd",x"c3",x"86"),
  2397 => (x"c3",x"87",x"d0",x"e5"),
  2398 => (x"ca",x"e5",x"49",x"fa"),
  2399 => (x"87",x"ce",x"c7",x"87"),
  2400 => (x"ff",x"c3",x"49",x"75"),
  2401 => (x"2d",x"b7",x"c8",x"99"),
  2402 => (x"9d",x"75",x"b5",x"71"),
  2403 => (x"87",x"e0",x"c0",x"02"),
  2404 => (x"7e",x"bf",x"c8",x"ff"),
  2405 => (x"dd",x"c2",x"49",x"6e"),
  2406 => (x"c2",x"89",x"bf",x"f4"),
  2407 => (x"c0",x"03",x"a9",x"e0"),
  2408 => (x"4d",x"c0",x"87",x"c5"),
  2409 => (x"c2",x"87",x"cf",x"c0"),
  2410 => (x"6e",x"48",x"f4",x"dd"),
  2411 => (x"87",x"c6",x"c0",x"78"),
  2412 => (x"48",x"f4",x"dd",x"c2"),
  2413 => (x"49",x"75",x"78",x"c0"),
  2414 => (x"c0",x"05",x"99",x"c8"),
  2415 => (x"f5",x"c3",x"87",x"ce"),
  2416 => (x"87",x"c3",x"e4",x"49"),
  2417 => (x"99",x"c2",x"49",x"70"),
  2418 => (x"87",x"ea",x"c0",x"02"),
  2419 => (x"bf",x"fc",x"f9",x"c2"),
  2420 => (x"87",x"ca",x"c0",x"02"),
  2421 => (x"c2",x"88",x"c1",x"48"),
  2422 => (x"c0",x"58",x"c0",x"fa"),
  2423 => (x"66",x"c4",x"87",x"d3"),
  2424 => (x"80",x"e0",x"c1",x"48"),
  2425 => (x"bf",x"6e",x"7e",x"70"),
  2426 => (x"87",x"c5",x"c0",x"02"),
  2427 => (x"73",x"49",x"ff",x"4b"),
  2428 => (x"48",x"a6",x"c8",x"0f"),
  2429 => (x"49",x"75",x"78",x"c1"),
  2430 => (x"c0",x"05",x"99",x"c4"),
  2431 => (x"f2",x"c3",x"87",x"ce"),
  2432 => (x"87",x"c3",x"e3",x"49"),
  2433 => (x"99",x"c2",x"49",x"70"),
  2434 => (x"87",x"f1",x"c0",x"02"),
  2435 => (x"bf",x"fc",x"f9",x"c2"),
  2436 => (x"c7",x"48",x"6e",x"7e"),
  2437 => (x"c0",x"03",x"a8",x"b7"),
  2438 => (x"48",x"6e",x"87",x"cb"),
  2439 => (x"fa",x"c2",x"80",x"c1"),
  2440 => (x"d3",x"c0",x"58",x"c0"),
  2441 => (x"48",x"66",x"c4",x"87"),
  2442 => (x"70",x"80",x"e0",x"c1"),
  2443 => (x"02",x"bf",x"6e",x"7e"),
  2444 => (x"4b",x"87",x"c5",x"c0"),
  2445 => (x"0f",x"73",x"49",x"fe"),
  2446 => (x"c1",x"48",x"a6",x"c8"),
  2447 => (x"49",x"fd",x"c3",x"78"),
  2448 => (x"70",x"87",x"c4",x"e2"),
  2449 => (x"02",x"99",x"c2",x"49"),
  2450 => (x"c2",x"87",x"e6",x"c0"),
  2451 => (x"02",x"bf",x"fc",x"f9"),
  2452 => (x"c2",x"87",x"c9",x"c0"),
  2453 => (x"c0",x"48",x"fc",x"f9"),
  2454 => (x"87",x"d0",x"c0",x"78"),
  2455 => (x"c1",x"4a",x"66",x"c4"),
  2456 => (x"02",x"6a",x"82",x"e0"),
  2457 => (x"4b",x"87",x"c5",x"c0"),
  2458 => (x"0f",x"73",x"49",x"fd"),
  2459 => (x"c1",x"48",x"a6",x"c8"),
  2460 => (x"49",x"fa",x"c3",x"78"),
  2461 => (x"70",x"87",x"d0",x"e1"),
  2462 => (x"02",x"99",x"c2",x"49"),
  2463 => (x"c2",x"87",x"ed",x"c0"),
  2464 => (x"48",x"bf",x"fc",x"f9"),
  2465 => (x"03",x"a8",x"b7",x"c7"),
  2466 => (x"c2",x"87",x"c9",x"c0"),
  2467 => (x"c7",x"48",x"fc",x"f9"),
  2468 => (x"87",x"d3",x"c0",x"78"),
  2469 => (x"c1",x"48",x"66",x"c4"),
  2470 => (x"7e",x"70",x"80",x"e0"),
  2471 => (x"c0",x"02",x"bf",x"6e"),
  2472 => (x"fc",x"4b",x"87",x"c5"),
  2473 => (x"c8",x"0f",x"73",x"49"),
  2474 => (x"78",x"c1",x"48",x"a6"),
  2475 => (x"f0",x"c3",x"48",x"75"),
  2476 => (x"48",x"7e",x"70",x"98"),
  2477 => (x"ce",x"c0",x"05",x"98"),
  2478 => (x"49",x"da",x"c1",x"87"),
  2479 => (x"70",x"87",x"c8",x"e0"),
  2480 => (x"02",x"99",x"c2",x"49"),
  2481 => (x"6e",x"87",x"ca",x"c1"),
  2482 => (x"87",x"cd",x"c0",x"05"),
  2483 => (x"ff",x"49",x"da",x"c1"),
  2484 => (x"70",x"87",x"f4",x"df"),
  2485 => (x"e8",x"c0",x"02",x"98"),
  2486 => (x"49",x"bf",x"e8",x"87"),
  2487 => (x"9b",x"ff",x"c3",x"4b"),
  2488 => (x"71",x"29",x"b7",x"c8"),
  2489 => (x"d9",x"db",x"ff",x"b3"),
  2490 => (x"c3",x"49",x"73",x"87"),
  2491 => (x"99",x"71",x"99",x"f0"),
  2492 => (x"87",x"e5",x"ff",x"05"),
  2493 => (x"ff",x"49",x"da",x"c1"),
  2494 => (x"70",x"87",x"cc",x"df"),
  2495 => (x"d8",x"ff",x"05",x"98"),
  2496 => (x"fc",x"f9",x"c2",x"87"),
  2497 => (x"cc",x"4b",x"49",x"bf"),
  2498 => (x"83",x"66",x"c4",x"93"),
  2499 => (x"73",x"71",x"4b",x"6b"),
  2500 => (x"02",x"9c",x"74",x"0f"),
  2501 => (x"6c",x"87",x"e9",x"c0"),
  2502 => (x"87",x"e4",x"c0",x"02"),
  2503 => (x"de",x"ff",x"49",x"6c"),
  2504 => (x"49",x"70",x"87",x"e5"),
  2505 => (x"c0",x"02",x"99",x"c1"),
  2506 => (x"a4",x"c4",x"87",x"cb"),
  2507 => (x"fc",x"f9",x"c2",x"4b"),
  2508 => (x"4b",x"6b",x"49",x"bf"),
  2509 => (x"02",x"84",x"c8",x"0f"),
  2510 => (x"6c",x"87",x"c5",x"c0"),
  2511 => (x"87",x"dc",x"ff",x"05"),
  2512 => (x"c0",x"02",x"66",x"c8"),
  2513 => (x"f9",x"c2",x"87",x"c8"),
  2514 => (x"f1",x"49",x"bf",x"fc"),
  2515 => (x"8e",x"ec",x"87",x"de"),
  2516 => (x"4c",x"26",x"4d",x"26"),
  2517 => (x"4f",x"26",x"4b",x"26"),
  2518 => (x"00",x"00",x"00",x"10"),
  2519 => (x"14",x"11",x"12",x"58"),
  2520 => (x"23",x"1c",x"1b",x"1d"),
  2521 => (x"94",x"91",x"59",x"5a"),
  2522 => (x"f4",x"eb",x"f2",x"f5"),
  2523 => (x"00",x"00",x"00",x"00"),
  2524 => (x"00",x"00",x"00",x"00"),
  2525 => (x"00",x"00",x"00",x"00"),
  2526 => (x"00",x"00",x"00",x"00"),
  2527 => (x"5c",x"5b",x"5e",x"0e"),
  2528 => (x"4b",x"71",x"0e",x"5d"),
  2529 => (x"d0",x"4c",x"d4",x"ff"),
  2530 => (x"78",x"c0",x"48",x"66"),
  2531 => (x"dd",x"ff",x"49",x"d6"),
  2532 => (x"ff",x"c3",x"87",x"f2"),
  2533 => (x"c3",x"49",x"6c",x"7c"),
  2534 => (x"4d",x"71",x"99",x"ff"),
  2535 => (x"99",x"f0",x"c3",x"49"),
  2536 => (x"05",x"a9",x"e0",x"c1"),
  2537 => (x"ff",x"c3",x"87",x"cb"),
  2538 => (x"c3",x"48",x"6c",x"7c"),
  2539 => (x"08",x"66",x"d0",x"98"),
  2540 => (x"7c",x"ff",x"c3",x"78"),
  2541 => (x"c8",x"49",x"4a",x"6c"),
  2542 => (x"7c",x"ff",x"c3",x"31"),
  2543 => (x"b2",x"71",x"4a",x"6c"),
  2544 => (x"31",x"c8",x"49",x"72"),
  2545 => (x"6c",x"7c",x"ff",x"c3"),
  2546 => (x"72",x"b2",x"71",x"4a"),
  2547 => (x"c3",x"31",x"c8",x"49"),
  2548 => (x"4a",x"6c",x"7c",x"ff"),
  2549 => (x"d0",x"ff",x"b2",x"71"),
  2550 => (x"78",x"e0",x"c0",x"48"),
  2551 => (x"c2",x"02",x"9b",x"73"),
  2552 => (x"75",x"7b",x"72",x"87"),
  2553 => (x"26",x"4d",x"26",x"48"),
  2554 => (x"26",x"4b",x"26",x"4c"),
  2555 => (x"4f",x"26",x"1e",x"4f"),
  2556 => (x"5c",x"5b",x"5e",x"0e"),
  2557 => (x"76",x"86",x"f8",x"0e"),
  2558 => (x"49",x"a6",x"c8",x"1e"),
  2559 => (x"c4",x"87",x"fd",x"fd"),
  2560 => (x"6e",x"4b",x"70",x"86"),
  2561 => (x"01",x"a8",x"c3",x"48"),
  2562 => (x"73",x"87",x"f4",x"c2"),
  2563 => (x"9a",x"f0",x"c3",x"4a"),
  2564 => (x"02",x"aa",x"d0",x"c1"),
  2565 => (x"e0",x"c1",x"87",x"c7"),
  2566 => (x"e2",x"c2",x"05",x"aa"),
  2567 => (x"c8",x"49",x"73",x"87"),
  2568 => (x"87",x"c3",x"02",x"99"),
  2569 => (x"73",x"87",x"c6",x"ff"),
  2570 => (x"c2",x"9c",x"c3",x"4c"),
  2571 => (x"c4",x"c1",x"05",x"ac"),
  2572 => (x"49",x"66",x"c4",x"87"),
  2573 => (x"1e",x"71",x"31",x"c9"),
  2574 => (x"c1",x"4a",x"66",x"c4"),
  2575 => (x"fa",x"c2",x"92",x"cc"),
  2576 => (x"81",x"72",x"49",x"c4"),
  2577 => (x"87",x"e6",x"ce",x"fe"),
  2578 => (x"da",x"ff",x"49",x"d8"),
  2579 => (x"c0",x"c8",x"87",x"f6"),
  2580 => (x"fc",x"e6",x"c2",x"1e"),
  2581 => (x"fc",x"e7",x"fd",x"49"),
  2582 => (x"48",x"d0",x"ff",x"87"),
  2583 => (x"c2",x"78",x"e0",x"c0"),
  2584 => (x"cc",x"1e",x"fc",x"e6"),
  2585 => (x"cc",x"c1",x"4a",x"66"),
  2586 => (x"c4",x"fa",x"c2",x"92"),
  2587 => (x"fe",x"81",x"72",x"49"),
  2588 => (x"cc",x"87",x"fc",x"cc"),
  2589 => (x"05",x"ac",x"c1",x"86"),
  2590 => (x"c4",x"87",x"c4",x"c1"),
  2591 => (x"31",x"c9",x"49",x"66"),
  2592 => (x"66",x"c4",x"1e",x"71"),
  2593 => (x"92",x"cc",x"c1",x"4a"),
  2594 => (x"49",x"c4",x"fa",x"c2"),
  2595 => (x"cd",x"fe",x"81",x"72"),
  2596 => (x"e6",x"c2",x"87",x"dc"),
  2597 => (x"66",x"c8",x"1e",x"fc"),
  2598 => (x"92",x"cc",x"c1",x"4a"),
  2599 => (x"49",x"c4",x"fa",x"c2"),
  2600 => (x"cb",x"fe",x"81",x"72"),
  2601 => (x"49",x"d7",x"87",x"ca"),
  2602 => (x"87",x"d8",x"d9",x"ff"),
  2603 => (x"c2",x"1e",x"c0",x"c8"),
  2604 => (x"fd",x"49",x"fc",x"e6"),
  2605 => (x"cc",x"87",x"fb",x"e5"),
  2606 => (x"48",x"d0",x"ff",x"86"),
  2607 => (x"f8",x"78",x"e0",x"c0"),
  2608 => (x"26",x"4c",x"26",x"8e"),
  2609 => (x"1e",x"4f",x"26",x"4b"),
  2610 => (x"b7",x"c4",x"4a",x"71"),
  2611 => (x"87",x"ce",x"03",x"aa"),
  2612 => (x"cc",x"c1",x"49",x"72"),
  2613 => (x"c4",x"fa",x"c2",x"91"),
  2614 => (x"81",x"c8",x"c1",x"81"),
  2615 => (x"4f",x"26",x"79",x"c0"),
  2616 => (x"5c",x"5b",x"5e",x"0e"),
  2617 => (x"86",x"fc",x"0e",x"5d"),
  2618 => (x"d4",x"ff",x"4a",x"71"),
  2619 => (x"d4",x"4c",x"c0",x"4b"),
  2620 => (x"b7",x"c3",x"4d",x"66"),
  2621 => (x"c2",x"c2",x"01",x"ad"),
  2622 => (x"02",x"9a",x"72",x"87"),
  2623 => (x"1e",x"87",x"ec",x"c0"),
  2624 => (x"cc",x"c1",x"49",x"75"),
  2625 => (x"c4",x"fa",x"c2",x"91"),
  2626 => (x"c8",x"80",x"71",x"48"),
  2627 => (x"66",x"c4",x"58",x"a6"),
  2628 => (x"e7",x"c4",x"fe",x"49"),
  2629 => (x"70",x"86",x"c4",x"87"),
  2630 => (x"87",x"d4",x"02",x"98"),
  2631 => (x"c8",x"c1",x"49",x"6e"),
  2632 => (x"6e",x"79",x"c1",x"81"),
  2633 => (x"69",x"81",x"c8",x"49"),
  2634 => (x"75",x"87",x"c5",x"4c"),
  2635 => (x"87",x"d7",x"fe",x"49"),
  2636 => (x"c8",x"48",x"d0",x"ff"),
  2637 => (x"7b",x"dd",x"78",x"e1"),
  2638 => (x"ff",x"c3",x"48",x"74"),
  2639 => (x"74",x"7b",x"70",x"98"),
  2640 => (x"29",x"b7",x"c8",x"49"),
  2641 => (x"ff",x"c3",x"48",x"71"),
  2642 => (x"74",x"7b",x"70",x"98"),
  2643 => (x"29",x"b7",x"d0",x"49"),
  2644 => (x"ff",x"c3",x"48",x"71"),
  2645 => (x"74",x"7b",x"70",x"98"),
  2646 => (x"28",x"b7",x"d8",x"48"),
  2647 => (x"7b",x"c0",x"7b",x"70"),
  2648 => (x"7b",x"7b",x"7b",x"7b"),
  2649 => (x"7b",x"7b",x"7b",x"7b"),
  2650 => (x"ff",x"7b",x"7b",x"7b"),
  2651 => (x"e0",x"c0",x"48",x"d0"),
  2652 => (x"dc",x"1e",x"75",x"78"),
  2653 => (x"f0",x"d6",x"ff",x"49"),
  2654 => (x"fc",x"86",x"c4",x"87"),
  2655 => (x"26",x"4d",x"26",x"8e"),
  2656 => (x"26",x"4b",x"26",x"4c"),
  2657 => (x"00",x"1c",x"e7",x"4f"),
  2658 => (x"00",x"1c",x"e7",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

