library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity DIAG10 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of DIAG10 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"78",X"D8",X"A2",X"00",X"BD",X"6C",X"C8",X"9D",X"00",X"B5",X"9D",X"00",X"B7",X"9D",X"00",X"99",
		X"9D",X"00",X"9B",X"E8",X"D0",X"EE",X"A9",X"FF",X"95",X"00",X"9D",X"00",X"01",X"9D",X"00",X"A0",
		X"9D",X"00",X"A1",X"9D",X"00",X"A2",X"9D",X"00",X"A3",X"9D",X"00",X"A4",X"9D",X"00",X"A5",X"9D",
		X"00",X"A6",X"9D",X"00",X"A7",X"9D",X"00",X"A8",X"9D",X"00",X"A9",X"9D",X"00",X"AA",X"9D",X"00",
		X"AB",X"9D",X"00",X"AC",X"9D",X"00",X"AD",X"9D",X"00",X"AE",X"9D",X"00",X"AF",X"9D",X"00",X"B0",
		X"9D",X"00",X"B1",X"9D",X"00",X"B2",X"9D",X"00",X"B3",X"9D",X"00",X"B4",X"9D",X"00",X"B6",X"9D",
		X"00",X"B8",X"9D",X"00",X"B9",X"9D",X"00",X"BA",X"9D",X"00",X"BB",X"9D",X"00",X"BC",X"9D",X"00",
		X"BD",X"9D",X"00",X"BE",X"9D",X"00",X"BF",X"E8",X"D0",X"9E",X"35",X"00",X"3D",X"00",X"01",X"3D",
		X"00",X"A0",X"3D",X"00",X"A1",X"3D",X"00",X"A2",X"3D",X"00",X"A3",X"3D",X"00",X"A4",X"3D",X"00",
		X"A5",X"3D",X"00",X"A6",X"3D",X"00",X"A7",X"3D",X"00",X"A8",X"3D",X"00",X"A9",X"3D",X"00",X"AA",
		X"3D",X"00",X"AB",X"3D",X"00",X"AC",X"3D",X"00",X"AD",X"3D",X"00",X"AE",X"3D",X"00",X"AF",X"3D",
		X"00",X"B0",X"3D",X"00",X"B1",X"3D",X"00",X"B2",X"3D",X"00",X"B3",X"3D",X"00",X"B4",X"3D",X"00",
		X"B6",X"3D",X"00",X"B8",X"3D",X"00",X"B9",X"3D",X"00",X"BA",X"3D",X"00",X"BB",X"3D",X"00",X"BC",
		X"3D",X"00",X"BD",X"3D",X"00",X"BE",X"3D",X"00",X"BF",X"E8",X"D0",X"9E",X"A8",X"A9",X"00",X"95",
		X"00",X"9D",X"00",X"01",X"9D",X"00",X"A0",X"9D",X"00",X"A1",X"9D",X"00",X"A2",X"9D",X"00",X"A3",
		X"9D",X"00",X"A4",X"9D",X"00",X"A5",X"9D",X"00",X"A6",X"9D",X"00",X"A7",X"9D",X"00",X"A8",X"9D",
		X"00",X"A9",X"9D",X"00",X"AA",X"9D",X"00",X"AB",X"9D",X"00",X"AC",X"9D",X"00",X"AD",X"9D",X"00",
		X"AE",X"9D",X"00",X"AF",X"9D",X"00",X"B0",X"9D",X"00",X"B1",X"9D",X"00",X"B2",X"9D",X"00",X"B3",
		X"9D",X"00",X"B4",X"9D",X"00",X"B6",X"9D",X"00",X"B8",X"9D",X"00",X"B9",X"9D",X"00",X"BA",X"9D",
		X"00",X"BB",X"9D",X"00",X"BC",X"9D",X"00",X"BD",X"9D",X"00",X"BE",X"9D",X"00",X"BF",X"E8",X"D0",
		X"9E",X"15",X"00",X"1D",X"00",X"01",X"1D",X"00",X"A0",X"1D",X"00",X"A1",X"1D",X"00",X"A2",X"1D",
		X"00",X"A3",X"1D",X"00",X"A4",X"1D",X"00",X"A5",X"1D",X"00",X"A6",X"1D",X"00",X"A7",X"1D",X"00",
		X"A8",X"1D",X"00",X"A9",X"1D",X"00",X"AA",X"1D",X"00",X"AB",X"1D",X"00",X"AC",X"1D",X"00",X"AD",
		X"1D",X"00",X"AE",X"1D",X"00",X"AF",X"1D",X"00",X"B0",X"1D",X"00",X"B1",X"1D",X"00",X"B2",X"1D",
		X"00",X"B3",X"1D",X"00",X"B4",X"1D",X"00",X"B6",X"1D",X"00",X"B8",X"1D",X"00",X"B9",X"1D",X"00",
		X"BA",X"1D",X"00",X"BB",X"1D",X"00",X"BC",X"1D",X"00",X"BD",X"1D",X"00",X"BE",X"1D",X"00",X"BF",
		X"E8",X"D0",X"9E",X"AA",X"4C",X"01",X"C2",X"C0",X"FF",X"D0",X"07",X"E0",X"00",X"D0",X"03",X"4C",
		X"9F",X"C6",X"98",X"49",X"FF",X"29",X"3F",X"D0",X"2F",X"8A",X"29",X"3F",X"D0",X"2A",X"8A",X"0A",
		X"0A",X"B0",X"04",X"98",X"49",X"40",X"0A",X"8A",X"30",X"03",X"98",X"30",X"0D",X"A2",X"FF",X"E8",
		X"BD",X"1C",X"C8",X"9D",X"90",X"BF",X"D0",X"F7",X"90",X"0B",X"A2",X"FF",X"E8",X"BD",X"13",X"C8",
		X"9D",X"A4",X"BF",X"D0",X"F7",X"38",X"B0",X"FE",X"8A",X"30",X"16",X"98",X"10",X"13",X"8A",X"29",
		X"60",X"D0",X"0E",X"8A",X"29",X"10",X"D0",X"04",X"A9",X"80",X"D0",X"05",X"8A",X"29",X"08",X"F0",
		X"F7",X"8E",X"06",X"03",X"8C",X"07",X"03",X"A2",X"00",X"A9",X"20",X"18",X"9D",X"80",X"BB",X"69",
		X"01",X"E8",X"E0",X"60",X"D0",X"F6",X"A2",X"00",X"BD",X"6C",X"C9",X"9D",X"00",X"99",X"9D",X"00",
		X"B5",X"BD",X"6C",X"CA",X"9D",X"00",X"9A",X"9D",X"00",X"B6",X"BD",X"6C",X"CB",X"9D",X"00",X"9B",
		X"9D",X"00",X"B7",X"E8",X"D0",X"E2",X"A0",X"14",X"A9",X"7F",X"9D",X"68",X"BF",X"9D",X"90",X"BF",
		X"9D",X"B8",X"BF",X"E8",X"88",X"D0",X"F3",X"A9",X"A0",X"A0",X"14",X"E0",X"28",X"D0",X"EB",X"A9",
		X"FF",X"8D",X"03",X"03",X"A9",X"FF",X"8D",X"00",X"03",X"A9",X"F7",X"8D",X"02",X"03",X"A9",X"CC",
		X"8D",X"0C",X"03",X"A9",X"07",X"8D",X"01",X"03",X"A9",X"EE",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",
		X"0C",X"03",X"A9",X"FF",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",
		X"03",X"A9",X"08",X"8D",X"01",X"03",X"A9",X"EE",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",
		X"AD",X"07",X"03",X"49",X"FF",X"0D",X"06",X"03",X"8D",X"06",X"03",X"A2",X"00",X"BD",X"6C",X"CC",
		X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",
		X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"6C",X"CC",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",
		X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",X"D0",X"CD",
		X"BD",X"6C",X"CD",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",
		X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"6C",X"CD",X"29",X"0F",X"8D",X"01",
		X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",
		X"E8",X"D0",X"CD",X"CA",X"D0",X"FD",X"88",X"D0",X"FA",X"A0",X"19",X"A2",X"C3",X"AD",X"06",X"03",
		X"4A",X"90",X"03",X"4C",X"1C",X"C6",X"4C",X"99",X"C5",X"8D",X"06",X"03",X"BD",X"6C",X"CE",X"4A",
		X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",
		X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"6C",X"CE",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",
		X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",X"D0",X"CD",X"CA",
		X"D0",X"FD",X"88",X"D0",X"FA",X"A0",X"65",X"A2",X"C3",X"AD",X"06",X"03",X"4A",X"90",X"03",X"4C",
		X"1C",X"C6",X"4C",X"99",X"C5",X"8D",X"06",X"03",X"BD",X"6C",X"CF",X"4A",X"4A",X"4A",X"4A",X"8D",
		X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",
		X"FD",X"BD",X"6C",X"CF",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",
		X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",X"D0",X"CD",X"CA",X"D0",X"FD",X"88",X"D0",
		X"FA",X"A0",X"B1",X"A2",X"C3",X"AD",X"06",X"03",X"4A",X"90",X"03",X"4C",X"1C",X"C6",X"4C",X"99",
		X"C5",X"8D",X"06",X"03",X"BD",X"67",X"D0",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",
		X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"67",X"D0",
		X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",
		X"30",X"88",X"D0",X"FD",X"E8",X"D0",X"CD",X"BD",X"67",X"D1",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",
		X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",
		X"BD",X"67",X"D1",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",
		X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",X"D0",X"CD",X"CA",X"D0",X"FD",X"88",X"D0",X"FA",
		X"A0",X"30",X"A2",X"C4",X"AD",X"06",X"03",X"4A",X"90",X"03",X"4C",X"1C",X"C6",X"4C",X"99",X"C5",
		X"8D",X"06",X"03",X"BD",X"67",X"D2",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",
		X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"67",X"D2",X"29",
		X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",
		X"88",X"D0",X"FD",X"E8",X"D0",X"CD",X"CA",X"D0",X"FD",X"88",X"D0",X"FA",X"A0",X"7C",X"A2",X"C4",
		X"AD",X"06",X"03",X"4A",X"90",X"03",X"4C",X"1C",X"C6",X"4C",X"99",X"C5",X"8D",X"06",X"03",X"BD",
		X"67",X"D3",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",
		X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"67",X"D3",X"29",X"0F",X"8D",X"01",X"03",
		X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",
		X"D0",X"CD",X"BD",X"67",X"D4",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",
		X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"67",X"D4",X"29",X"0F",
		X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",
		X"D0",X"FD",X"E8",X"D0",X"CD",X"CA",X"D0",X"FD",X"88",X"D0",X"FA",X"A0",X"FB",X"A2",X"C4",X"AD",
		X"06",X"03",X"4A",X"90",X"03",X"4C",X"1C",X"C6",X"4C",X"99",X"C5",X"8D",X"06",X"03",X"BD",X"67",
		X"D5",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",
		X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"BD",X"67",X"D5",X"29",X"0F",X"8D",X"01",X"03",X"A9",
		X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",X"D0",
		X"CD",X"CA",X"D0",X"FD",X"88",X"D0",X"FA",X"A0",X"47",X"A2",X"C5",X"AD",X"06",X"03",X"4A",X"90",
		X"03",X"4C",X"1C",X"C6",X"4C",X"99",X"C5",X"8D",X"06",X"03",X"BD",X"67",X"D6",X"4A",X"4A",X"4A",
		X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",
		X"88",X"D0",X"FD",X"BD",X"67",X"D6",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",
		X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"30",X"88",X"D0",X"FD",X"E8",X"D0",X"CD",X"CA",X"D0",X"FD",
		X"88",X"D0",X"FA",X"A0",X"93",X"A2",X"C5",X"AD",X"06",X"03",X"4A",X"90",X"03",X"4C",X"1C",X"C6",
		X"4C",X"99",X"C5",X"8D",X"06",X"03",X"38",X"B0",X"FE",X"8C",X"06",X"03",X"8E",X"07",X"03",X"A8",
		X"A2",X"00",X"BD",X"62",X"D7",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",
		X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"38",X"A9",X"30",X"E9",X"01",X"D0",X"FC",X"BD",X"62",X"D7",
		X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"38",
		X"A9",X"30",X"E9",X"01",X"D0",X"FC",X"E8",X"D0",X"C9",X"BD",X"62",X"D8",X"4A",X"4A",X"4A",X"4A",
		X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"38",X"A9",X"30",
		X"E9",X"01",X"D0",X"FC",X"BD",X"62",X"D8",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",
		X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"38",X"A9",X"30",X"E9",X"01",X"D0",X"FC",X"E8",X"D0",X"C9",
		X"38",X"E9",X"01",X"D0",X"FB",X"CA",X"D0",X"F8",X"98",X"6C",X"06",X"03",X"8C",X"06",X"03",X"8E",
		X"07",X"03",X"A8",X"A2",X"00",X"BD",X"61",X"D9",X"4A",X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",
		X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"38",X"A9",X"30",X"E9",X"01",X"D0",X"FC",
		X"BD",X"61",X"D9",X"29",X"0F",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",
		X"0C",X"03",X"38",X"A9",X"30",X"E9",X"01",X"D0",X"FC",X"E8",X"D0",X"C9",X"BD",X"61",X"DA",X"4A",
		X"4A",X"4A",X"4A",X"8D",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",
		X"38",X"A9",X"30",X"E9",X"01",X"D0",X"FC",X"BD",X"61",X"DA",X"29",X"0F",X"8D",X"01",X"03",X"A9",
		X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"38",X"A9",X"30",X"E9",X"01",X"D0",X"FC",
		X"E8",X"D0",X"C9",X"38",X"E9",X"01",X"D0",X"FB",X"CA",X"D0",X"F8",X"98",X"6C",X"06",X"03",X"20",
		X"8A",X"C7",X"A9",X"C8",X"A0",X"25",X"20",X"C1",X"C7",X"20",X"C4",X"C7",X"A9",X"C8",X"A0",X"3C",
		X"20",X"C1",X"C7",X"A9",X"FF",X"8D",X"03",X"03",X"A9",X"FF",X"8D",X"00",X"03",X"A9",X"F7",X"8D",
		X"02",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A9",X"7F",X"8D",X"0D",X"03",X"AD",X"0D",X"03",X"D0",
		X"20",X"A9",X"0A",X"8D",X"06",X"03",X"A9",X"00",X"8D",X"05",X"03",X"AD",X"04",X"03",X"C9",X"06",
		X"D0",X"0F",X"AD",X"0D",X"03",X"F0",X"0A",X"A9",X"C8",X"A0",X"43",X"20",X"C1",X"C7",X"4C",X"FB",
		X"C6",X"A9",X"C8",X"A0",X"4B",X"20",X"C1",X"C7",X"38",X"B0",X"FE",X"A9",X"07",X"A2",X"FE",X"20",
		X"D5",X"C7",X"A9",X"00",X"A2",X"18",X"20",X"D5",X"C7",X"A9",X"01",X"A2",X"00",X"20",X"D5",X"C7",
		X"A9",X"08",X"A2",X"10",X"20",X"D5",X"C7",X"A9",X"0C",X"A2",X"0F",X"20",X"D5",X"C7",X"A9",X"00",
		X"20",X"F0",X"C7",X"E0",X"18",X"F0",X"0A",X"A9",X"C8",X"A0",X"5B",X"20",X"C1",X"C7",X"38",X"B0",
		X"FE",X"A9",X"C8",X"A0",X"54",X"20",X"C1",X"C7",X"20",X"C4",X"C7",X"A9",X"C8",X"A0",X"63",X"20",
		X"C1",X"C7",X"A9",X"0E",X"8D",X"01",X"03",X"A9",X"EE",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",
		X"03",X"A9",X"60",X"85",X"12",X"A9",X"BD",X"85",X"13",X"A9",X"FE",X"48",X"8D",X"01",X"03",X"A9",
		X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A0",X"07",X"98",X"09",X"F8",X"8D",X"00",
		X"03",X"A9",X"08",X"2C",X"00",X"03",X"F0",X"02",X"09",X"80",X"91",X"12",X"88",X"10",X"EC",X"20",
		X"C4",X"C7",X"68",X"38",X"2A",X"B0",X"D4",X"4C",X"51",X"C7",X"A9",X"1A",X"8D",X"DF",X"BF",X"A9",
		X"80",X"85",X"12",X"A9",X"BB",X"85",X"13",X"A9",X"00",X"8D",X"67",X"02",X"60",X"84",X"10",X"85",
		X"11",X"A0",X"00",X"B1",X"10",X"F0",X"19",X"E6",X"10",X"D0",X"02",X"E6",X"11",X"AC",X"67",X"02",
		X"91",X"12",X"C8",X"8C",X"67",X"02",X"C0",X"28",X"D0",X"E7",X"20",X"C4",X"C7",X"4C",X"A1",X"C7",
		X"60",X"20",X"9D",X"C7",X"18",X"A5",X"12",X"69",X"28",X"85",X"12",X"90",X"02",X"E6",X"13",X"A9",
		X"00",X"8D",X"67",X"02",X"60",X"8D",X"01",X"03",X"A9",X"EE",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",
		X"0C",X"03",X"8E",X"01",X"03",X"A9",X"EC",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"60",
		X"8D",X"01",X"03",X"A9",X"EE",X"8D",X"0C",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"A9",X"CE",X"8D",
		X"0C",X"03",X"AE",X"01",X"03",X"A9",X"CC",X"8D",X"0C",X"03",X"60",X"01",X"02",X"04",X"08",X"10",
		X"20",X"40",X"80",X"62",X"61",X"64",X"20",X"69",X"63",X"79",X"7C",X"00",X"62",X"61",X"64",X"20",
		X"69",X"63",X"79",X"7D",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"72",X"6F",X"6D",X"20",X"64",X"69",X"61",X"67",X"20",X"77",X"00",X"72",X"61",X"6D",X"20",
		X"6F",X"6B",X"00",X"7C",X"7B",X"78",X"78",X"20",X"6F",X"6B",X"00",X"62",X"61",X"64",X"20",X"7C",
		X"7B",X"78",X"78",X"00",X"70",X"73",X"67",X"20",X"6F",X"6B",X"00",X"62",X"61",X"64",X"20",X"70",
		X"73",X"67",X"00",X"6B",X"62",X"64",X"20",X"74",X"65",X"73",X"74",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"14",X"22",X"22",X"3E",X"22",X"22",X"00",X"3C",X"22",X"22",X"3C",
		X"22",X"22",X"3C",X"00",X"1C",X"22",X"20",X"20",X"20",X"22",X"1C",X"00",X"3C",X"22",X"22",X"22",
		X"22",X"22",X"3C",X"00",X"3E",X"20",X"20",X"3C",X"20",X"20",X"3E",X"00",X"3E",X"20",X"20",X"3C",
		X"20",X"20",X"20",X"00",X"1E",X"20",X"20",X"20",X"26",X"22",X"1E",X"00",X"22",X"22",X"22",X"3E",
		X"22",X"22",X"22",X"00",X"1C",X"08",X"08",X"08",X"08",X"08",X"1C",X"00",X"02",X"02",X"02",X"02",
		X"02",X"22",X"1C",X"00",X"22",X"24",X"28",X"30",X"28",X"24",X"22",X"00",X"20",X"20",X"20",X"20",
		X"20",X"20",X"3E",X"00",X"22",X"36",X"2A",X"2A",X"22",X"22",X"22",X"00",X"22",X"22",X"32",X"2A",
		X"26",X"22",X"22",X"00",X"1C",X"22",X"22",X"22",X"22",X"22",X"1C",X"00",X"3C",X"22",X"22",X"3C",
		X"20",X"20",X"20",X"00",X"1C",X"22",X"22",X"22",X"2A",X"24",X"1A",X"00",X"3C",X"22",X"22",X"3C",
		X"28",X"24",X"22",X"00",X"1C",X"22",X"20",X"1C",X"02",X"22",X"1C",X"00",X"3E",X"08",X"08",X"08",
		X"08",X"08",X"08",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"1C",X"00",X"1C",X"22",X"26",X"2A",
		X"32",X"22",X"1C",X"00",X"08",X"18",X"08",X"08",X"08",X"08",X"1C",X"00",X"1C",X"22",X"02",X"04",
		X"08",X"10",X"3E",X"00",X"3E",X"02",X"04",X"0C",X"02",X"22",X"1C",X"00",X"04",X"0C",X"14",X"24",
		X"3E",X"04",X"04",X"00",X"3E",X"20",X"3C",X"02",X"02",X"22",X"1C",X"00",X"0C",X"10",X"20",X"3C",
		X"22",X"22",X"1C",X"00",X"3E",X"02",X"04",X"08",X"10",X"10",X"10",X"00",X"1C",X"22",X"22",X"1C",
		X"22",X"22",X"1C",X"00",X"1C",X"22",X"22",X"1E",X"02",X"04",X"18",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"33",X"2D",X"2D",X"2D",X"33",X"3F",X"3F",X"3F",X"37",X"27",X"37",
		X"37",X"23",X"3F",X"3F",X"3F",X"37",X"27",X"37",X"37",X"23",X"3F",X"00",X"3F",X"0F",X"37",X"2F",
		X"1F",X"07",X"3F",X"3F",X"3F",X"0F",X"37",X"2F",X"1F",X"07",X"3F",X"00",X"3F",X"0F",X"37",X"2F",
		X"1F",X"07",X"3F",X"00",X"3F",X"0F",X"37",X"2F",X"1F",X"07",X"3F",X"00",X"3F",X"39",X"3E",X"3D",
		X"3E",X"39",X"3F",X"3F",X"3F",X"0F",X"2F",X"0F",X"2F",X"0F",X"3F",X"00",X"3F",X"0F",X"2F",X"0F",
		X"2F",X"0F",X"3F",X"00",X"3F",X"0F",X"2F",X"0F",X"2F",X"0F",X"3F",X"00",X"3F",X"0F",X"2F",X"0F",
		X"2F",X"0F",X"3F",X"00",X"3F",X"0F",X"2F",X"0F",X"2F",X"0F",X"3F",X"00",X"3F",X"0F",X"2F",X"0F",
		X"2F",X"0F",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"37",X"35",X"31",
		X"3D",X"3D",X"3F",X"3F",X"3F",X"37",X"35",X"31",X"3D",X"3D",X"3F",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3D",X"1D",X"1C",
		X"1F",X"1F",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3D",X"1D",X"1C",
		X"1F",X"1F",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3D",X"1D",X"1C",
		X"1F",X"1F",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"10",X"1C",X"14",X"1C",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"06",X"01",X"06",X"00",X"3F",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"06",X"01",X"06",X"00",X"3F",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"10",X"18",X"04",X"18",X"00",X"00",X"00",X"1C",X"10",X"18",
		X"04",X"18",X"00",X"3F",X"00",X"1C",X"10",X"18",X"04",X"18",X"00",X"00",X"3F",X"33",X"2F",X"23",
		X"2B",X"23",X"3F",X"3F",X"3F",X"33",X"2F",X"23",X"2B",X"23",X"3F",X"00",X"3F",X"33",X"2F",X"23",
		X"2B",X"23",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"27",X"1F",X"07",
		X"17",X"07",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"23",X"20",X"20",X"00",X"3F",X"3F",X"3C",X"3B",X"38",
		X"3A",X"38",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"23",X"20",X"20",X"00",X"3F",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"0E",
		X"02",X"02",X"00",X"3F",X"00",X"08",X"0A",X"0E",X"02",X"02",X"00",X"00",X"3F",X"3C",X"3B",X"38",
		X"3A",X"38",X"3F",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"30",X"10",X"30",X"00",X"3F",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"30",X"10",X"30",X"00",X"3F",X"00",X"30",X"10",X"30",
		X"10",X"30",X"00",X"3F",X"00",X"06",X"01",X"02",X"01",X"06",X"00",X"00",X"07",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"08",X"10",X"20",X"38",X"00",X"3F",X"00",X"30",X"08",X"10",
		X"20",X"38",X"00",X"3F",X"00",X"30",X"08",X"10",X"20",X"38",X"00",X"00",X"00",X"08",X"18",X"08",
		X"08",X"1C",X"00",X"3F",X"00",X"08",X"18",X"08",X"08",X"1C",X"00",X"00",X"00",X"0C",X"12",X"12",
		X"12",X"0C",X"00",X"00",X"07",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"98",X"88",
		X"87",X"88",X"89",X"89",X"88",X"88",X"88",X"78",X"77",X"77",X"77",X"78",X"89",X"99",X"99",X"98",
		X"87",X"77",X"88",X"89",X"98",X"88",X"88",X"77",X"77",X"77",X"77",X"77",X"78",X"99",X"AA",X"99",
		X"88",X"77",X"77",X"89",X"99",X"99",X"88",X"87",X"87",X"88",X"88",X"77",X"77",X"67",X"79",X"9A",
		X"AA",X"99",X"87",X"77",X"78",X"99",X"A9",X"98",X"77",X"77",X"88",X"87",X"77",X"66",X"67",X"8A",
		X"AB",X"AA",X"97",X"76",X"77",X"8A",X"AA",X"A8",X"87",X"87",X"78",X"88",X"77",X"65",X"57",X"7A",
		X"BB",X"C9",X"A8",X"67",X"57",X"89",X"AA",X"A8",X"97",X"88",X"78",X"78",X"76",X"65",X"53",X"97",
		X"DC",X"CC",X"99",X"66",X"57",X"89",X"B9",X"B8",X"88",X"78",X"78",X"78",X"76",X"54",X"54",X"89",
		X"CC",X"CA",X"97",X"67",X"69",X"9B",X"BA",X"97",X"87",X"88",X"88",X"77",X"65",X"54",X"49",X"8D",
		X"CB",X"C7",X"75",X"57",X"7A",X"AB",X"A9",X"87",X"88",X"88",X"88",X"76",X"55",X"54",X"69",X"AD",
		X"CC",X"A8",X"76",X"67",X"8A",X"AA",X"A8",X"88",X"89",X"88",X"87",X"76",X"66",X"66",X"59",X"9B",
		X"CA",X"A8",X"77",X"67",X"88",X"9A",X"99",X"98",X"88",X"88",X"77",X"77",X"77",X"77",X"77",X"78",
		X"99",X"B9",X"99",X"77",X"77",X"88",X"99",X"99",X"88",X"88",X"87",X"77",X"78",X"88",X"88",X"87",
		X"77",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"87",X"77",X"77",X"89",X"99",X"99",X"88",X"88",X"87",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"87",X"77",X"77",X"77",X"89",X"A9",X"99",X"88",X"77",X"88",X"88",X"99",X"98",X"88",X"88",
		X"88",X"88",X"87",X"77",X"77",X"77",X"78",X"AB",X"A9",X"88",X"87",X"77",X"89",X"99",X"98",X"88",
		X"88",X"88",X"77",X"77",X"77",X"77",X"76",X"68",X"AB",X"A9",X"88",X"88",X"77",X"89",X"AA",X"98",
		X"88",X"88",X"88",X"88",X"87",X"77",X"66",X"66",X"8A",X"BB",X"A9",X"88",X"77",X"78",X"9A",X"A9",
		X"98",X"88",X"88",X"88",X"88",X"77",X"66",X"65",X"68",X"BC",X"B9",X"88",X"87",X"67",X"89",X"AA",
		X"98",X"88",X"88",X"88",X"87",X"77",X"66",X"65",X"68",X"AC",X"BA",X"98",X"87",X"66",X"79",X"AA",
		X"A9",X"88",X"88",X"88",X"87",X"77",X"77",X"66",X"67",X"8A",X"BB",X"99",X"88",X"77",X"67",X"89",
		X"A9",X"99",X"88",X"88",X"87",X"77",X"77",X"77",X"76",X"78",X"9A",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"99",
		X"99",X"88",X"88",X"87",X"77",X"77",X"77",X"77",X"7B",X"B9",X"98",X"8A",X"98",X"78",X"99",X"89",
		X"88",X"87",X"87",X"77",X"77",X"77",X"66",X"8B",X"A9",X"88",X"9A",X"88",X"88",X"99",X"88",X"88",
		X"87",X"87",X"77",X"77",X"66",X"66",X"8B",X"AA",X"98",X"AA",X"88",X"88",X"98",X"88",X"88",X"78",
		X"87",X"77",X"77",X"66",X"66",X"67",X"CB",X"A9",X"89",X"B9",X"98",X"69",X"89",X"97",X"87",X"78",
		X"77",X"77",X"76",X"77",X"66",X"57",X"DC",X"A9",X"79",X"B9",X"98",X"89",X"88",X"88",X"87",X"88",
		X"77",X"77",X"76",X"55",X"44",X"CF",X"CB",X"98",X"A9",X"88",X"68",X"98",X"98",X"89",X"88",X"87",
		X"88",X"77",X"75",X"55",X"55",X"4D",X"FB",X"B9",X"8B",X"98",X"86",X"8A",X"98",X"78",X"99",X"87",
		X"78",X"87",X"65",X"54",X"56",X"5A",X"FC",X"CA",X"8A",X"98",X"87",X"89",X"98",X"88",X"99",X"97",
		X"78",X"77",X"76",X"65",X"56",X"76",X"9D",X"BB",X"A8",X"99",X"88",X"77",X"88",X"99",X"89",X"99",
		X"87",X"77",X"77",X"76",X"65",X"66",X"65",X"CB",X"BA",X"99",X"A9",X"87",X"78",X"89",X"A9",X"98",
		X"88",X"87",X"77",X"87",X"76",X"66",X"66",X"57",X"BB",X"BA",X"9A",X"A8",X"87",X"78",X"99",X"98",
		X"98",X"88",X"77",X"78",X"88",X"77",X"66",X"66",X"65",X"9C",X"BB",X"99",X"A9",X"87",X"78",X"99",
		X"98",X"88",X"88",X"87",X"88",X"88",X"87",X"66",X"66",X"65",X"8B",X"BB",X"99",X"99",X"88",X"78",
		X"89",X"98",X"88",X"88",X"87",X"78",X"88",X"87",X"76",X"66",X"66",X"7A",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"88",X"87",
		X"78",X"88",X"88",X"88",X"87",X"77",X"77",X"78",X"89",X"99",X"99",X"99",X"99",X"99",X"98",X"88",
		X"87",X"77",X"77",X"66",X"55",X"47",X"79",X"AB",X"DC",X"CA",X"87",X"55",X"66",X"9A",X"BB",X"BA",
		X"87",X"65",X"55",X"54",X"33",X"68",X"CD",X"DF",X"DC",X"96",X"54",X"56",X"8B",X"CD",X"CB",X"97",
		X"64",X"44",X"44",X"32",X"77",X"AD",X"EF",X"EB",X"A7",X"55",X"36",X"9A",X"CC",X"CB",X"98",X"65",
		X"54",X"44",X"31",X"66",X"AD",X"FF",X"FC",X"B8",X"54",X"25",X"8A",X"DD",X"DC",X"98",X"65",X"54",
		X"43",X"21",X"67",X"BD",X"EF",X"EC",X"A7",X"54",X"35",X"89",X"CC",X"CB",X"98",X"65",X"54",X"43",
		X"12",X"57",X"DE",X"EF",X"DC",X"96",X"54",X"36",X"7A",X"DC",X"CA",X"98",X"65",X"55",X"43",X"12",
		X"57",X"CE",X"EF",X"DC",X"96",X"54",X"46",X"7A",X"CC",X"CA",X"98",X"66",X"65",X"54",X"21",X"56",
		X"AC",X"EF",X"FC",X"A8",X"55",X"34",X"68",X"AC",X"CC",X"A9",X"87",X"66",X"54",X"32",X"15",X"7B",
		X"DE",X"FE",X"DA",X"86",X"53",X"46",X"9B",X"BC",X"CB",X"A8",X"76",X"55",X"33",X"21",X"57",X"CE",
		X"EF",X"FD",X"B7",X"54",X"24",X"57",X"AB",X"CC",X"CB",X"97",X"65",X"44",X"33",X"25",X"6A",X"DF",
		X"FF",X"CB",X"85",X"43",X"35",X"7A",X"CC",X"DC",X"B9",X"76",X"54",X"44",X"33",X"37",X"7A",X"DE",
		X"FF",X"CB",X"75",X"42",X"45",X"7A",X"BD",X"DC",X"C9",X"86",X"44",X"44",X"55",X"56",X"69",X"9C",
		X"CC",X"CB",X"A8",X"65",X"55",X"67",X"9A",X"BC",X"BB",X"98",X"75",X"55",X"56",X"67",X"87",X"77",
		X"88",X"9A",X"AA",X"AA",X"98",X"77",X"77",X"79",X"9A",X"AA",X"98",X"76",X"66",X"77",X"89",X"99",
		X"87",X"65",X"56",X"78",X"AA",X"BB",X"BA",X"99",X"87",X"9A",X"97",X"78",X"88",X"87",X"88",X"88",
		X"77",X"88",X"88",X"78",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"98",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"78",
		X"87",X"77",X"88",X"88",X"88",X"98",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"99",X"98",X"77",X"88",X"99",X"88",X"88",X"88",X"88",X"88",X"87",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"87",X"88",X"88",X"99",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"88",X"77",
		X"78",X"99",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"78",X"88",X"88",
		X"77",X"77",X"89",X"AA",X"A9",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"77",X"77",
		X"77",X"77",X"76",X"68",X"AC",X"BA",X"87",X"78",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"87",
		X"77",X"77",X"77",X"65",X"57",X"AD",X"DB",X"86",X"68",X"99",X"88",X"89",X"99",X"98",X"78",X"88",
		X"87",X"77",X"77",X"77",X"75",X"57",X"BE",X"EA",X"65",X"79",X"A9",X"87",X"89",X"AA",X"87",X"77",
		X"88",X"77",X"67",X"77",X"76",X"53",X"6B",X"FF",X"A5",X"36",X"BC",X"A7",X"57",X"9B",X"A8",X"67",
		X"89",X"98",X"77",X"78",X"87",X"66",X"55",X"8D",X"FC",X"74",X"6A",X"CA",X"75",X"79",X"AA",X"87",
		X"78",X"98",X"77",X"78",X"77",X"65",X"53",X"6C",X"FF",X"72",X"4B",X"EB",X"64",X"6A",X"BA",X"87",
		X"79",X"98",X"77",X"88",X"77",X"66",X"64",X"39",X"FF",X"A2",X"2A",X"FD",X"74",X"6A",X"BA",X"87",
		X"79",X"98",X"77",X"87",X"66",X"66",X"53",X"4B",X"FF",X"62",X"7E",X"E9",X"45",X"8A",X"BB",X"96",
		X"79",X"A9",X"87",X"76",X"66",X"65",X"32",X"9F",X"F7",X"27",X"DD",X"84",X"58",X"9A",X"A8",X"67",
		X"9A",X"98",X"87",X"76",X"66",X"54",X"26",X"EF",X"B3",X"4B",X"FB",X"65",X"78",X"9A",X"97",X"79",
		X"A9",X"87",X"88",X"76",X"55",X"54",X"39",X"FF",X"73",X"8D",X"C8",X"66",X"78",X"AA",X"86",X"7A",
		X"B9",X"77",X"78",X"76",X"65",X"54",X"4A",X"FC",X"65",X"AC",X"A8",X"67",X"79",X"A9",X"77",X"8A",
		X"A8",X"78",X"87",X"76",X"76",X"66",X"58",X"CC",X"86",X"8A",X"A9",X"87",X"78",X"99",X"88",X"99",
		X"88",X"88",X"87",X"66",X"77",X"77",X"76",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"A9",X"A7",X"98",X"88",X"89",X"88",X"88",X"87",X"88",
		X"78",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"89",X"98",X"88",X"87",X"76",X"54",X"48",X"8F",
		X"BE",X"99",X"57",X"8B",X"BB",X"89",X"67",X"44",X"10",X"0C",X"AF",X"CE",X"35",X"48",X"CC",X"F8",
		X"B4",X"A6",X"A8",X"84",X"00",X"0F",X"CF",X"AB",X"01",X"8C",X"FD",X"A3",X"59",X"AC",X"88",X"54",
		X"20",X"02",X"FE",X"F2",X"40",X"6F",X"FE",X"60",X"7A",X"FC",X"64",X"5A",X"55",X"10",X"1F",X"FF",
		X"40",X"17",X"FF",X"95",X"07",X"FF",X"E0",X"58",X"BA",X"64",X"00",X"3F",X"FF",X"00",X"4F",X"FF",
		X"10",X"0D",X"FE",X"60",X"7D",X"B8",X"72",X"00",X"3F",X"FF",X"00",X"7F",X"FF",X"00",X"3F",X"F8",
		X"32",X"BE",X"A8",X"71",X"00",X"1F",X"FF",X"00",X"6F",X"FF",X"00",X"6F",X"FB",X"05",X"AD",X"A6",
		X"82",X"00",X"1F",X"FB",X"10",X"3F",X"FE",X"00",X"5F",X"FB",X"04",X"AC",X"A8",X"95",X"00",X"1F",
		X"FD",X"40",X"1F",X"FE",X"30",X"0F",X"FC",X"22",X"9C",X"B9",X"A6",X"00",X"17",X"FF",X"30",X"1F",
		X"FF",X"30",X"1F",X"FF",X"22",X"6C",X"E9",X"A7",X"11",X"11",X"FF",X"71",X"15",X"FF",X"61",X"17",
		X"FF",X"31",X"4B",X"FB",X"87",X"51",X"11",X"BF",X"F1",X"11",X"EF",X"F1",X"11",X"BF",X"F2",X"19",
		X"CF",X"96",X"73",X"11",X"2F",X"FC",X"12",X"4F",X"FD",X"11",X"4D",X"FF",X"11",X"9E",X"F9",X"47",
		X"41",X"13",X"FF",X"C3",X"14",X"FF",X"E5",X"02",X"8F",X"F9",X"44",X"AE",X"C7",X"56",X"40",X"1B",
		X"FF",X"A8",X"45",X"BD",X"CA",X"85",X"57",X"AB",X"A9",X"77",X"8A",X"A9",X"76",X"77",X"88",X"88",
		X"88",X"8A",X"AA",X"87",X"79",X"A9",X"86",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"87",X"66",X"54",X"43",
		X"79",X"BD",X"BB",X"A9",X"A9",X"9A",X"9C",X"BA",X"A9",X"99",X"88",X"78",X"88",X"87",X"75",X"43",
		X"21",X"2A",X"BD",X"B7",X"87",X"9A",X"88",X"78",X"99",X"A9",X"88",X"78",X"88",X"88",X"88",X"76",
		X"53",X"32",X"3A",X"EE",X"D8",X"AB",X"CC",X"87",X"67",X"AC",X"B9",X"89",X"9A",X"87",X"77",X"98",
		X"64",X"32",X"11",X"07",X"EC",X"E7",X"AC",X"BD",X"77",X"77",X"B8",X"86",X"69",X"89",X"88",X"9A",
		X"BA",X"88",X"67",X"55",X"43",X"20",X"37",X"EB",X"B8",X"AC",X"CB",X"78",X"78",X"A7",X"87",X"9A",
		X"B9",X"98",X"AA",X"99",X"77",X"65",X"54",X"31",X"01",X"CC",X"DB",X"6D",X"AD",X"A6",X"87",X"AA",
		X"A8",X"89",X"9A",X"78",X"79",X"A9",X"87",X"87",X"77",X"56",X"43",X"22",X"3E",X"AD",X"AA",X"CC",
		X"B7",X"86",X"9A",X"89",X"A9",X"B9",X"98",X"88",X"89",X"88",X"77",X"76",X"65",X"53",X"22",X"4D",
		X"AE",X"99",X"CB",X"B8",X"86",X"99",X"99",X"89",X"99",X"87",X"88",X"99",X"88",X"87",X"77",X"77",
		X"65",X"43",X"23",X"99",X"DB",X"8C",X"AC",X"98",X"69",X"89",X"9A",X"9A",X"99",X"88",X"88",X"98",
		X"98",X"77",X"77",X"65",X"54",X"42",X"39",X"9D",X"BA",X"BC",X"CA",X"97",X"98",X"98",X"87",X"88",
		X"98",X"88",X"9A",X"A9",X"88",X"88",X"77",X"66",X"54",X"43",X"33",X"A8",X"CA",X"BB",X"DA",X"B8",
		X"88",X"98",X"88",X"98",X"A9",X"88",X"98",X"A9",X"98",X"88",X"87",X"77",X"76",X"54",X"42",X"35",
		X"7C",X"AB",X"CC",X"BB",X"98",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"89",X"88",X"87",X"77",
		X"76",X"65",X"44",X"43",X"56",X"BB",X"BC",X"BB",X"B9",X"88",X"78",X"88",X"89",X"AA",X"99",X"9A",
		X"A9",X"88",X"77",X"77",X"66",X"65",X"54",X"43",X"5C",X"8B",X"CA",X"CB",X"A9",X"87",X"78",X"88",
		X"89",X"99",X"98",X"99",X"99",X"88",X"88",X"77",X"77",X"76",X"66",X"55",X"44",X"69",X"9A",X"AA",
		X"BB",X"A9",X"88",X"88",X"88",X"89",X"99",X"99",X"99",X"99",X"88",X"88",X"87",X"77",X"77",X"76",
		X"65",X"55",X"68",X"99",X"AA",X"AA",X"A9",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"77",X"77",X"66",X"55",X"56",X"78",X"9A",X"AA",X"AA",X"99",X"88",X"88",X"88",X"88",
		X"89",X"88",X"88",X"88",X"88",X"88",X"87",X"77",X"76",X"65",X"55",X"67",X"89",X"AA",X"AA",X"A9",
		X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"87",X"77",X"66",X"65",
		X"56",X"78",X"9A",X"AA",X"AA",X"A9",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"77",X"66",X"66",X"66",X"78",X"9A",X"AA",X"AA",X"99",X"98",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"77",X"66",X"66",X"67",X"89",X"9A",X"AA",X"A9",X"99",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"77",X"76",X"66",X"67",X"89",
		X"9A",X"AA",X"A9",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"77",X"76",X"67",X"78",X"9A",X"BB",X"BA",X"99",X"87",
		X"77",X"77",X"78",X"88",X"88",X"77",X"66",X"66",X"78",X"9A",X"BB",X"BB",X"A9",X"87",X"77",X"78",
		X"89",X"99",X"88",X"77",X"66",X"55",X"55",X"78",X"AB",X"CC",X"CA",X"97",X"76",X"76",X"88",X"99",
		X"99",X"98",X"77",X"66",X"55",X"54",X"68",X"AB",X"CC",X"CB",X"A8",X"76",X"66",X"78",X"99",X"9A",
		X"99",X"87",X"66",X"54",X"44",X"67",X"AB",X"CC",X"CB",X"A8",X"86",X"76",X"77",X"88",X"99",X"99",
		X"88",X"76",X"55",X"54",X"56",X"9A",X"CC",X"CC",X"B9",X"87",X"66",X"67",X"78",X"9A",X"A9",X"98",
		X"76",X"44",X"45",X"69",X"AB",X"BC",X"CC",X"A9",X"77",X"66",X"67",X"89",X"9A",X"A9",X"98",X"75",
		X"54",X"45",X"69",X"AB",X"BC",X"CC",X"A9",X"77",X"66",X"67",X"78",X"9A",X"A9",X"98",X"76",X"54",
		X"45",X"68",X"9A",X"AC",X"CC",X"AA",X"87",X"66",X"56",X"78",X"9A",X"AA",X"99",X"86",X"54",X"45",
		X"68",X"89",X"AB",X"CC",X"BA",X"98",X"66",X"56",X"78",X"9A",X"AA",X"A9",X"87",X"65",X"55",X"66",
		X"79",X"AC",X"CC",X"BA",X"98",X"66",X"56",X"68",X"89",X"AA",X"A9",X"87",X"75",X"54",X"56",X"88",
		X"AA",X"BB",X"BA",X"A8",X"86",X"66",X"77",X"89",X"9A",X"A9",X"98",X"77",X"65",X"55",X"67",X"89",
		X"AB",X"BB",X"A9",X"87",X"76",X"67",X"78",X"99",X"99",X"98",X"87",X"77",X"66",X"67",X"78",X"89",
		X"AA",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"9A",X"AA",X"99",X"98",X"88",X"77",X"77",X"65",X"55",
		X"44",X"99",X"EC",X"CB",X"89",X"79",X"8A",X"99",X"98",X"87",X"88",X"87",X"76",X"54",X"32",X"2C",
		X"BF",X"DA",X"95",X"88",X"9A",X"A9",X"89",X"7A",X"89",X"88",X"76",X"75",X"52",X"20",X"C8",X"FF",
		X"9C",X"29",X"7A",X"C8",X"A6",X"97",X"AA",X"89",X"79",X"79",X"67",X"54",X"21",X"0B",X"9F",X"F9",
		X"B2",X"98",X"BC",X"99",X"58",X"7C",X"BA",X"87",X"A8",X"A6",X"74",X"52",X"00",X"9A",X"FF",X"9C",
		X"29",X"8A",X"D9",X"95",X"77",X"99",X"9A",X"8A",X"89",X"77",X"66",X"54",X"31",X"1C",X"AF",X"DB",
		X"86",X"77",X"B8",X"A7",X"77",X"7A",X"BC",X"A9",X"88",X"87",X"76",X"65",X"43",X"27",X"9E",X"FB",
		X"D6",X"86",X"79",X"8A",X"89",X"79",X"99",X"A9",X"98",X"87",X"76",X"77",X"77",X"66",X"57",X"8A",
		X"CB",X"B9",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"87",X"77",X"76",X"65",X"56",X"8A",
		X"AB",X"AA",X"AA",X"98",X"76",X"67",X"89",X"AA",X"A9",X"98",X"87",X"65",X"55",X"55",X"57",X"9B",
		X"CC",X"BA",X"A9",X"98",X"66",X"67",X"89",X"AA",X"AA",X"98",X"86",X"65",X"55",X"54",X"57",X"9B",
		X"CC",X"BB",X"AA",X"98",X"65",X"56",X"89",X"AA",X"AA",X"98",X"87",X"66",X"55",X"54",X"56",X"8A",
		X"BC",X"CB",X"BA",X"A9",X"76",X"55",X"68",X"9A",X"AA",X"98",X"88",X"87",X"65",X"55",X"55",X"57",
		X"9B",X"CC",X"CB",X"AA",X"98",X"65",X"67",X"9A",X"AA",X"98",X"89",X"87",X"65",X"55",X"54",X"46",
		X"8B",X"CC",X"CB",X"BA",X"98",X"65",X"56",X"89",X"A9",X"99",X"99",X"87",X"66",X"55",X"43",X"35",
		X"8A",X"CC",X"CB",X"BB",X"97",X"54",X"57",X"89",X"99",X"99",X"88",X"76",X"67",X"76",X"53",X"35",
		X"8A",X"CE",X"FF",X"FD",X"A6",X"55",X"78",X"9A",X"BC",X"CA",X"98",X"87",X"65",X"43",X"22",X"47",
		X"AB",X"BC",X"DC",X"96",X"44",X"32",X"47",X"9B",X"CC",X"CC",X"BA",X"86",X"53",X"10",X"14",X"7A",
		X"DF",X"FF",X"B8",X"76",X"54",X"69",X"BC",X"DF",X"FD",X"A8",X"64",X"32",X"10",X"04",X"8A",X"DF",
		X"FF",X"ED",X"96",X"44",X"34",X"8A",X"BD",X"ED",X"A9",X"52",X"00",X"00",X"01",X"38",X"FF",X"FF",
		X"FC",X"97",X"21",X"01",X"58",X"AC",X"DD",X"DC",X"86",X"51",X"00",X"25",X"AF",X"FF",X"FF",X"FF",
		X"A7",X"31",X"33",X"69",X"BD",X"DD",X"B8",X"62",X"00",X"00",X"01",X"7B",X"EF",X"FF",X"EC",X"94",
		X"41",X"24",X"6A",X"AD",X"DC",X"B7",X"63",X"10",X"03",X"18",X"7D",X"FF",X"FF",X"FB",X"B8",X"48",
		X"48",X"98",X"DA",X"DC",X"99",X"43",X"00",X"30",X"44",X"6F",X"AF",X"CE",X"D8",X"A4",X"65",X"45",
		X"67",X"9B",X"AB",X"96",X"52",X"13",X"02",X"67",X"DD",X"FE",X"EC",X"BB",X"88",X"56",X"56",X"88",
		X"AA",X"A9",X"76",X"43",X"30",X"26",X"9B",X"CE",X"CE",X"DD",X"C9",X"97",X"65",X"67",X"89",X"A9",
		X"98",X"75",X"42",X"46",X"44",X"5A",X"CE",X"ED",X"C9",X"A8",X"88",X"77",X"67",X"78",X"99",X"97",
		X"65",X"32",X"27",X"89",X"78",X"AC",X"FD",X"DA",X"98",X"77",X"56",X"78",X"98",X"99",X"88",X"65",
		X"33",X"26",X"8A",X"88",X"AC",X"EE",X"DB",X"98",X"77",X"66",X"77",X"99",X"99",X"98",X"75",X"43",
		X"36",X"77",X"68",X"AD",X"ED",X"CA",X"A9",X"77",X"67",X"67",X"88",X"AA",X"99",X"76",X"54",X"43",
		X"34",X"7B",X"CD",X"CC",X"DC",X"C9",X"86",X"56",X"67",X"89",X"99",X"A9",X"87",X"64",X"34",X"55",
		X"66",X"9B",X"DE",X"DC",X"BA",X"98",X"65",X"66",X"78",X"99",X"AA",X"98",X"76",X"43",X"35",X"67",
		X"79",X"BD",X"ED",X"CA",X"98",X"77",X"66",X"67",X"89",X"AA",X"98",X"76",X"54",X"54",X"45",X"7A",
		X"BC",X"CC",X"CB",X"B9",X"86",X"56",X"78",X"88",X"99",X"99",X"87",X"65",X"44",X"56",X"78",X"9A",
		X"BC",X"CB",X"A9",X"98",X"76",X"77",X"88",X"89",X"99",X"88",X"76",X"55",X"55",X"67",X"89",X"AB",
		X"BB",X"BA",X"98",X"87",X"77",X"77",X"88",X"88",X"88",X"87",X"76",X"66",X"67",X"88",X"9A",X"AB",
		X"BB",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"99",X"99",X"99",X"98",X"88",X"77",X"76",X"66",X"56",X"78",X"99",X"AA",X"AA",X"AA",X"A9",
		X"99",X"98",X"88",X"77",X"76",X"66",X"55",X"66",X"78",X"9A",X"AA",X"AA",X"AA",X"99",X"99",X"88",
		X"88",X"87",X"77",X"77",X"65",X"55",X"67",X"89",X"AA",X"AB",X"AA",X"A9",X"98",X"88",X"88",X"88",
		X"88",X"87",X"76",X"65",X"44",X"56",X"79",X"9A",X"AB",X"BB",X"AA",X"98",X"88",X"88",X"88",X"88",
		X"88",X"77",X"66",X"54",X"45",X"67",X"9A",X"BB",X"BB",X"BA",X"A9",X"88",X"88",X"88",X"88",X"88",
		X"77",X"76",X"65",X"43",X"55",X"78",X"9B",X"BB",X"CB",X"BA",X"A9",X"99",X"88",X"88",X"87",X"77",
		X"77",X"76",X"54",X"34",X"56",X"89",X"BB",X"CC",X"CB",X"BA",X"99",X"99",X"88",X"88",X"77",X"77",
		X"77",X"66",X"54",X"34",X"57",X"9A",X"BC",X"CC",X"BB",X"AA",X"99",X"88",X"88",X"88",X"87",X"77",
		X"76",X"65",X"43",X"34",X"67",X"9B",X"BC",X"CC",X"BB",X"A9",X"89",X"88",X"88",X"88",X"88",X"77",
		X"76",X"65",X"43",X"34",X"67",X"9B",X"CC",X"CC",X"CB",X"AA",X"99",X"88",X"88",X"87",X"77",X"77",
		X"76",X"65",X"43",X"44",X"68",X"9B",X"BC",X"CC",X"BB",X"A9",X"98",X"98",X"88",X"88",X"87",X"77",
		X"76",X"54",X"32",X"44",X"68",X"AC",X"CC",X"DC",X"CB",X"A9",X"88",X"88",X"88",X"88",X"87",X"87",
		X"76",X"65",X"43",X"23",X"57",X"AB",X"CC",X"CC",X"CB",X"A9",X"89",X"88",X"88",X"88",X"88",X"77",
		X"77",X"65",X"44",X"24",X"47",X"8A",X"CC",X"DC",X"CC",X"AA",X"98",X"88",X"88",X"88",X"88",X"88",
		X"77",X"66",X"54",X"32",X"44",X"79",X"BC",X"CC",X"CC",X"BA",X"99",X"88",X"88",X"88",X"88",X"88",
		X"87",X"77",X"64",X"53",X"14",X"47",X"9B",X"CC",X"CC",X"CB",X"AA",X"99",X"99",X"98",X"98",X"77",
		X"77",X"66",X"30",X"00",X"18",X"BF",X"EA",X"BB",X"AD",X"96",X"83",X"7D",X"AC",X"A7",X"A9",X"8A",
		X"88",X"72",X"00",X"00",X"08",X"EF",X"FF",X"BF",X"BB",X"B5",X"14",X"7D",X"FB",X"79",X"9A",X"C9",
		X"79",X"50",X"00",X"00",X"4F",X"FF",X"E7",X"6F",X"F8",X"94",X"07",X"FD",X"A9",X"67",X"DD",X"99",
		X"85",X"10",X"00",X"01",X"FF",X"BC",X"B4",X"FF",X"B2",X"35",X"4E",X"F9",X"36",X"BA",X"CD",X"75",
		X"73",X"00",X"00",X"3F",X"F9",X"6D",X"BA",X"FF",X"20",X"5C",X"ED",X"A6",X"59",X"EB",X"87",X"76",
		X"10",X"00",X"0D",X"FF",X"46",X"DF",X"CC",X"B3",X"04",X"FF",X"A2",X"4A",X"CB",X"99",X"77",X"51",
		X"00",X"00",X"FF",X"D3",X"6F",X"FE",X"86",X"54",X"6E",X"FA",X"14",X"BF",X"B7",X"79",X"73",X"00",
		X"00",X"9F",X"F9",X"27",X"FF",X"D4",X"36",X"AB",X"DC",X"84",X"5A",X"DB",X"75",X"65",X"20",X"00",
		X"8F",X"FA",X"46",X"EF",X"F6",X"24",X"9E",X"DA",X"65",X"7A",X"B9",X"77",X"75",X"30",X"00",X"7F",
		X"FB",X"45",X"CF",X"F9",X"21",X"8F",X"FB",X"43",X"7B",X"C9",X"65",X"77",X"51",X"00",X"3D",X"FE",
		X"73",X"7F",X"FF",X"71",X"3A",X"FF",X"A3",X"26",X"CD",X"A6",X"45",X"65",X"20",X"04",X"DF",X"E8",
		X"58",X"EF",X"E7",X"33",X"8E",X"FA",X"52",X"59",X"CC",X"85",X"34",X"54",X"21",X"39",X"DE",X"C9",
		X"9B",X"DD",X"B8",X"67",X"9B",X"A8",X"66",X"68",X"99",X"86",X"43",X"33",X"56",X"9B",X"BB",X"AB",
		X"CB",X"A9",X"88",X"89",X"99",X"87",X"77",X"89",X"98",X"76",X"54",X"44",X"46",X"79",X"AB",X"BB",
		X"BA",X"9A",X"99",X"99",X"88",X"88",X"88",X"87",X"77",X"77",X"65",X"54",X"46",X"89",X"AB",X"BA",
		X"AA",X"A9",X"99",X"99",X"88",X"88",X"88",X"77",X"77",X"87",X"76",X"55",X"66",X"78",X"99",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
