
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"f9",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"c0",x"f9",x"c2"),
    14 => (x"48",x"cc",x"e6",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c7",x"e0"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"cc",x"e6"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"e6",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"cc"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"d0",x"e6",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"d4",x"e6",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"d4",x"e6"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"e6",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"d4"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"e6",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"db"),
   285 => (x"e6",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"dc"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"dd",x"e6",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"dd",x"e6",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"de",x"e6"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"e6",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"d9"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"da",x"e6"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"db",x"e6",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"dc",x"e6"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"fa",x"ee",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"f2",x"e6"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"cb",x"f2",x"c0"),
   331 => (x"e8",x"e7",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f2",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"c7"),
   337 => (x"71",x"4a",x"c4",x"e8"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"f8",x"ed",x"c2",x"87"),
   343 => (x"ee",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"f0"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"f8",x"ed",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"f2",x"e6",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f2",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"c7"),
   359 => (x"71",x"4a",x"c4",x"e8"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"ee",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"fa"),
   364 => (x"f2",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"cb"),
   366 => (x"71",x"4a",x"e8",x"e7"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"f0",x"ee",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"f1",x"ee",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"f2",x"e6"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"fd",x"e6"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"e6",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"fe"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"ff",x"e6"),
   394 => (x"f6",x"ee",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"ee",x"c2",x"88",x"c1"),
   397 => (x"e7",x"c2",x"58",x"fa"),
   398 => (x"49",x"bf",x"97",x"c0"),
   399 => (x"e7",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"c1"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"c7",x"f3",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"c2",x"e7"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"fa",x"ee",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"c7",x"f2",x"c0"),
   409 => (x"c4",x"e8",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"ee",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"f2"),
   416 => (x"c2",x"5c",x"db",x"f3"),
   417 => (x"bf",x"97",x"d7",x"e7"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"d6",x"e7"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"d8",x"e7"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"e7",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"d9"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"c7",x"f3",x"c2"),
   428 => (x"cf",x"f3",x"c2",x"81"),
   429 => (x"df",x"e7",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"de",x"e7",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"e0",x"e7",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"e1",x"e7",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"d3",x"f3",x"c2",x"4a"),
   440 => (x"cf",x"f3",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"f3",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"d3"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"c4",x"e7",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"c3",x"e7",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"c2",x"ef",x"c2"),
   450 => (x"bf",x"fe",x"ee",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"db",x"f3",x"c2"),
   454 => (x"97",x"c9",x"e7",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"c8",x"e7",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"d7",x"f3",x"c2",x"82"),
   460 => (x"cf",x"f3",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"cb",x"f3"),
   463 => (x"f3",x"c2",x"78",x"a1"),
   464 => (x"f3",x"c2",x"48",x"db"),
   465 => (x"c2",x"78",x"bf",x"cf"),
   466 => (x"c2",x"48",x"df",x"f3"),
   467 => (x"78",x"bf",x"d3",x"f3"),
   468 => (x"bf",x"fa",x"ee",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"d7",x"f3",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"ee",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"fe"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"fa",x"ee",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"c7",x"f3"),
   489 => (x"bf",x"c3",x"f2",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"c7",x"f2",x"c0"),
   492 => (x"1e",x"f2",x"e6",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"fa",x"ee",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"f2",x"e6",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"e6",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"f2"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"ca",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"ee"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"c2",x"ef"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"c9",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"ee"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"1e",x"0e",x"5d",x"5c"),
   533 => (x"05",x"9b",x"4b",x"71"),
   534 => (x"48",x"c0",x"87",x"c5"),
   535 => (x"c8",x"87",x"e5",x"c1"),
   536 => (x"7d",x"c0",x"4d",x"a3"),
   537 => (x"c7",x"02",x"66",x"d4"),
   538 => (x"97",x"66",x"d4",x"87"),
   539 => (x"87",x"c5",x"05",x"bf"),
   540 => (x"cf",x"c1",x"48",x"c0"),
   541 => (x"49",x"66",x"d4",x"87"),
   542 => (x"70",x"87",x"f3",x"fd"),
   543 => (x"c1",x"02",x"9c",x"4c"),
   544 => (x"a4",x"dc",x"87",x"c0"),
   545 => (x"da",x"7d",x"69",x"49"),
   546 => (x"a3",x"c4",x"49",x"a4"),
   547 => (x"7a",x"69",x"9f",x"4a"),
   548 => (x"bf",x"fa",x"ee",x"c2"),
   549 => (x"d4",x"87",x"d2",x"02"),
   550 => (x"69",x"9f",x"49",x"a4"),
   551 => (x"ff",x"ff",x"c0",x"49"),
   552 => (x"d0",x"48",x"71",x"99"),
   553 => (x"c2",x"7e",x"70",x"30"),
   554 => (x"6e",x"7e",x"c0",x"87"),
   555 => (x"80",x"6a",x"48",x"49"),
   556 => (x"7b",x"c0",x"7a",x"70"),
   557 => (x"6a",x"49",x"a3",x"cc"),
   558 => (x"49",x"a3",x"d0",x"79"),
   559 => (x"48",x"74",x"79",x"c0"),
   560 => (x"48",x"c0",x"87",x"c2"),
   561 => (x"87",x"ec",x"fa",x"26"),
   562 => (x"5c",x"5b",x"5e",x"0e"),
   563 => (x"4c",x"71",x"0e",x"5d"),
   564 => (x"48",x"c3",x"f2",x"c0"),
   565 => (x"9c",x"74",x"78",x"ff"),
   566 => (x"87",x"ca",x"c1",x"02"),
   567 => (x"69",x"49",x"a4",x"c8"),
   568 => (x"87",x"c2",x"c1",x"02"),
   569 => (x"6c",x"4a",x"66",x"d0"),
   570 => (x"a6",x"d4",x"82",x"49"),
   571 => (x"4d",x"66",x"d0",x"5a"),
   572 => (x"f6",x"ee",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e4",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"f4",x"f9",x"49"),
   578 => (x"ee",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"f2"),
   580 => (x"75",x"7c",x"71",x"81"),
   581 => (x"f6",x"ee",x"c2",x"b9"),
   582 => (x"ba",x"ff",x"4a",x"bf"),
   583 => (x"99",x"71",x"99",x"72"),
   584 => (x"87",x"dc",x"ff",x"05"),
   585 => (x"cb",x"f9",x"7c",x"75"),
   586 => (x"1e",x"73",x"1e",x"87"),
   587 => (x"02",x"9b",x"4b",x"71"),
   588 => (x"a3",x"c8",x"87",x"c7"),
   589 => (x"c5",x"05",x"69",x"49"),
   590 => (x"c0",x"48",x"c0",x"87"),
   591 => (x"f3",x"c2",x"87",x"eb"),
   592 => (x"c4",x"4a",x"bf",x"cb"),
   593 => (x"49",x"69",x"49",x"a3"),
   594 => (x"ee",x"c2",x"89",x"c2"),
   595 => (x"71",x"91",x"bf",x"f2"),
   596 => (x"ee",x"c2",x"4a",x"a2"),
   597 => (x"6b",x"49",x"bf",x"f6"),
   598 => (x"4a",x"a2",x"71",x"99"),
   599 => (x"72",x"1e",x"66",x"c8"),
   600 => (x"87",x"d2",x"ea",x"49"),
   601 => (x"49",x"70",x"86",x"c4"),
   602 => (x"87",x"cc",x"f8",x"48"),
   603 => (x"71",x"1e",x"73",x"1e"),
   604 => (x"c7",x"02",x"9b",x"4b"),
   605 => (x"49",x"a3",x"c8",x"87"),
   606 => (x"87",x"c5",x"05",x"69"),
   607 => (x"eb",x"c0",x"48",x"c0"),
   608 => (x"cb",x"f3",x"c2",x"87"),
   609 => (x"a3",x"c4",x"4a",x"bf"),
   610 => (x"c2",x"49",x"69",x"49"),
   611 => (x"f2",x"ee",x"c2",x"89"),
   612 => (x"a2",x"71",x"91",x"bf"),
   613 => (x"f6",x"ee",x"c2",x"4a"),
   614 => (x"99",x"6b",x"49",x"bf"),
   615 => (x"c8",x"4a",x"a2",x"71"),
   616 => (x"49",x"72",x"1e",x"66"),
   617 => (x"c4",x"87",x"c5",x"e6"),
   618 => (x"48",x"49",x"70",x"86"),
   619 => (x"0e",x"87",x"c9",x"f7"),
   620 => (x"5d",x"5c",x"5b",x"5e"),
   621 => (x"4b",x"71",x"1e",x"0e"),
   622 => (x"c9",x"4c",x"66",x"d4"),
   623 => (x"02",x"9b",x"73",x"2c"),
   624 => (x"c8",x"87",x"cf",x"c1"),
   625 => (x"02",x"69",x"49",x"a3"),
   626 => (x"d0",x"87",x"c7",x"c1"),
   627 => (x"66",x"d4",x"4d",x"a3"),
   628 => (x"f6",x"ee",x"c2",x"7d"),
   629 => (x"b9",x"ff",x"49",x"bf"),
   630 => (x"7e",x"99",x"4a",x"6b"),
   631 => (x"cd",x"03",x"ac",x"71"),
   632 => (x"7d",x"7b",x"c0",x"87"),
   633 => (x"c4",x"4a",x"a3",x"cc"),
   634 => (x"79",x"6a",x"49",x"a3"),
   635 => (x"8c",x"72",x"87",x"c2"),
   636 => (x"dd",x"02",x"9c",x"74"),
   637 => (x"73",x"1e",x"49",x"87"),
   638 => (x"87",x"cc",x"fb",x"49"),
   639 => (x"66",x"d4",x"86",x"c4"),
   640 => (x"99",x"ff",x"c7",x"49"),
   641 => (x"c2",x"87",x"cb",x"02"),
   642 => (x"73",x"1e",x"f2",x"e6"),
   643 => (x"87",x"d9",x"fc",x"49"),
   644 => (x"f5",x"26",x"86",x"c4"),
   645 => (x"73",x"1e",x"87",x"de"),
   646 => (x"9b",x"4b",x"71",x"1e"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"5b",x"df",x"f3",x"c2"),
   649 => (x"8a",x"c2",x"4a",x"73"),
   650 => (x"bf",x"f2",x"ee",x"c2"),
   651 => (x"f3",x"c2",x"92",x"49"),
   652 => (x"72",x"48",x"bf",x"cb"),
   653 => (x"e3",x"f3",x"c2",x"80"),
   654 => (x"c4",x"48",x"71",x"58"),
   655 => (x"c2",x"ef",x"c2",x"30"),
   656 => (x"87",x"ed",x"c0",x"58"),
   657 => (x"48",x"db",x"f3",x"c2"),
   658 => (x"bf",x"cf",x"f3",x"c2"),
   659 => (x"df",x"f3",x"c2",x"78"),
   660 => (x"d3",x"f3",x"c2",x"48"),
   661 => (x"ee",x"c2",x"78",x"bf"),
   662 => (x"c9",x"02",x"bf",x"fa"),
   663 => (x"f2",x"ee",x"c2",x"87"),
   664 => (x"31",x"c4",x"49",x"bf"),
   665 => (x"f3",x"c2",x"87",x"c7"),
   666 => (x"c4",x"49",x"bf",x"d7"),
   667 => (x"c2",x"ef",x"c2",x"31"),
   668 => (x"87",x"c4",x"f4",x"59"),
   669 => (x"5c",x"5b",x"5e",x"0e"),
   670 => (x"c0",x"4a",x"71",x"0e"),
   671 => (x"02",x"9a",x"72",x"4b"),
   672 => (x"da",x"87",x"e1",x"c0"),
   673 => (x"69",x"9f",x"49",x"a2"),
   674 => (x"fa",x"ee",x"c2",x"4b"),
   675 => (x"87",x"cf",x"02",x"bf"),
   676 => (x"9f",x"49",x"a2",x"d4"),
   677 => (x"c0",x"4c",x"49",x"69"),
   678 => (x"d0",x"9c",x"ff",x"ff"),
   679 => (x"c0",x"87",x"c2",x"34"),
   680 => (x"b3",x"49",x"74",x"4c"),
   681 => (x"ed",x"fd",x"49",x"73"),
   682 => (x"87",x"ca",x"f3",x"87"),
   683 => (x"5c",x"5b",x"5e",x"0e"),
   684 => (x"86",x"f4",x"0e",x"5d"),
   685 => (x"7e",x"c0",x"4a",x"71"),
   686 => (x"d8",x"02",x"9a",x"72"),
   687 => (x"ee",x"e6",x"c2",x"87"),
   688 => (x"c2",x"78",x"c0",x"48"),
   689 => (x"c2",x"48",x"e6",x"e6"),
   690 => (x"78",x"bf",x"df",x"f3"),
   691 => (x"48",x"ea",x"e6",x"c2"),
   692 => (x"bf",x"db",x"f3",x"c2"),
   693 => (x"cf",x"ef",x"c2",x"78"),
   694 => (x"c2",x"50",x"c0",x"48"),
   695 => (x"49",x"bf",x"fe",x"ee"),
   696 => (x"bf",x"ee",x"e6",x"c2"),
   697 => (x"03",x"aa",x"71",x"4a"),
   698 => (x"72",x"87",x"ff",x"c3"),
   699 => (x"05",x"99",x"cf",x"49"),
   700 => (x"c2",x"87",x"e0",x"c0"),
   701 => (x"c2",x"1e",x"f2",x"e6"),
   702 => (x"49",x"bf",x"e6",x"e6"),
   703 => (x"48",x"e6",x"e6",x"c2"),
   704 => (x"71",x"78",x"a1",x"c1"),
   705 => (x"c4",x"87",x"ef",x"e3"),
   706 => (x"ff",x"f1",x"c0",x"86"),
   707 => (x"f2",x"e6",x"c2",x"48"),
   708 => (x"c0",x"87",x"cc",x"78"),
   709 => (x"48",x"bf",x"ff",x"f1"),
   710 => (x"c0",x"80",x"e0",x"c0"),
   711 => (x"c2",x"58",x"c3",x"f2"),
   712 => (x"48",x"bf",x"ee",x"e6"),
   713 => (x"e6",x"c2",x"80",x"c1"),
   714 => (x"7f",x"27",x"58",x"f2"),
   715 => (x"bf",x"00",x"00",x"0c"),
   716 => (x"9d",x"4d",x"bf",x"97"),
   717 => (x"87",x"e2",x"c2",x"02"),
   718 => (x"02",x"ad",x"e5",x"c3"),
   719 => (x"c0",x"87",x"db",x"c2"),
   720 => (x"4b",x"bf",x"ff",x"f1"),
   721 => (x"11",x"49",x"a3",x"cb"),
   722 => (x"05",x"ac",x"cf",x"4c"),
   723 => (x"75",x"87",x"d2",x"c1"),
   724 => (x"c1",x"99",x"df",x"49"),
   725 => (x"c2",x"91",x"cd",x"89"),
   726 => (x"c1",x"81",x"c2",x"ef"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c3"),
   729 => (x"4a",x"a3",x"c5",x"51"),
   730 => (x"a3",x"c7",x"51",x"12"),
   731 => (x"c9",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"ce"),
   734 => (x"4a",x"a3",x"d0",x"51"),
   735 => (x"a3",x"d2",x"51",x"12"),
   736 => (x"d4",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"d6"),
   739 => (x"4a",x"a3",x"d8",x"51"),
   740 => (x"a3",x"dc",x"51",x"12"),
   741 => (x"de",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"f9",x"c0",x"7e",x"c1"),
   744 => (x"c8",x"49",x"74",x"87"),
   745 => (x"ea",x"c0",x"05",x"99"),
   746 => (x"d0",x"49",x"74",x"87"),
   747 => (x"87",x"d0",x"05",x"99"),
   748 => (x"c0",x"02",x"66",x"dc"),
   749 => (x"49",x"73",x"87",x"ca"),
   750 => (x"70",x"0f",x"66",x"dc"),
   751 => (x"87",x"d3",x"02",x"98"),
   752 => (x"c6",x"c0",x"05",x"6e"),
   753 => (x"c2",x"ef",x"c2",x"87"),
   754 => (x"c0",x"50",x"c0",x"48"),
   755 => (x"48",x"bf",x"ff",x"f1"),
   756 => (x"c2",x"87",x"e7",x"c2"),
   757 => (x"c0",x"48",x"cf",x"ef"),
   758 => (x"ee",x"c2",x"7e",x"50"),
   759 => (x"c2",x"49",x"bf",x"fe"),
   760 => (x"4a",x"bf",x"ee",x"e6"),
   761 => (x"fc",x"04",x"aa",x"71"),
   762 => (x"f3",x"c2",x"87",x"c1"),
   763 => (x"c0",x"05",x"bf",x"df"),
   764 => (x"ee",x"c2",x"87",x"c8"),
   765 => (x"c1",x"02",x"bf",x"fa"),
   766 => (x"f2",x"c0",x"87",x"fe"),
   767 => (x"78",x"ff",x"48",x"c3"),
   768 => (x"bf",x"ea",x"e6",x"c2"),
   769 => (x"87",x"f4",x"ed",x"49"),
   770 => (x"e6",x"c2",x"49",x"70"),
   771 => (x"a6",x"c4",x"59",x"ee"),
   772 => (x"ea",x"e6",x"c2",x"48"),
   773 => (x"ee",x"c2",x"78",x"bf"),
   774 => (x"c0",x"02",x"bf",x"fa"),
   775 => (x"66",x"c4",x"87",x"d8"),
   776 => (x"ff",x"ff",x"cf",x"49"),
   777 => (x"a9",x"99",x"f8",x"ff"),
   778 => (x"87",x"c5",x"c0",x"02"),
   779 => (x"e1",x"c0",x"4d",x"c0"),
   780 => (x"c0",x"4d",x"c1",x"87"),
   781 => (x"66",x"c4",x"87",x"dc"),
   782 => (x"f8",x"ff",x"cf",x"49"),
   783 => (x"c0",x"02",x"a9",x"99"),
   784 => (x"a6",x"c8",x"87",x"c8"),
   785 => (x"c0",x"78",x"c0",x"48"),
   786 => (x"a6",x"c8",x"87",x"c5"),
   787 => (x"c8",x"78",x"c1",x"48"),
   788 => (x"9d",x"75",x"4d",x"66"),
   789 => (x"87",x"e0",x"c0",x"05"),
   790 => (x"c2",x"49",x"66",x"c4"),
   791 => (x"f2",x"ee",x"c2",x"89"),
   792 => (x"c2",x"91",x"4a",x"bf"),
   793 => (x"4a",x"bf",x"cb",x"f3"),
   794 => (x"48",x"e6",x"e6",x"c2"),
   795 => (x"c2",x"78",x"a1",x"72"),
   796 => (x"c0",x"48",x"ee",x"e6"),
   797 => (x"87",x"e3",x"f9",x"78"),
   798 => (x"8e",x"f4",x"48",x"c0"),
   799 => (x"00",x"87",x"f5",x"eb"),
   800 => (x"ff",x"00",x"00",x"00"),
   801 => (x"8f",x"ff",x"ff",x"ff"),
   802 => (x"98",x"00",x"00",x"0c"),
   803 => (x"46",x"00",x"00",x"0c"),
   804 => (x"32",x"33",x"54",x"41"),
   805 => (x"00",x"20",x"20",x"20"),
   806 => (x"31",x"54",x"41",x"46"),
   807 => (x"20",x"20",x"20",x"36"),
   808 => (x"d4",x"ff",x"1e",x"00"),
   809 => (x"78",x"ff",x"c3",x"48"),
   810 => (x"4f",x"26",x"48",x"68"),
   811 => (x"48",x"d4",x"ff",x"1e"),
   812 => (x"ff",x"78",x"ff",x"c3"),
   813 => (x"e1",x"c8",x"48",x"d0"),
   814 => (x"48",x"d4",x"ff",x"78"),
   815 => (x"f3",x"c2",x"78",x"d4"),
   816 => (x"d4",x"ff",x"48",x"e3"),
   817 => (x"4f",x"26",x"50",x"bf"),
   818 => (x"48",x"d0",x"ff",x"1e"),
   819 => (x"26",x"78",x"e0",x"c0"),
   820 => (x"cc",x"ff",x"1e",x"4f"),
   821 => (x"99",x"49",x"70",x"87"),
   822 => (x"c0",x"87",x"c6",x"02"),
   823 => (x"f1",x"05",x"a9",x"fb"),
   824 => (x"26",x"48",x"71",x"87"),
   825 => (x"5b",x"5e",x"0e",x"4f"),
   826 => (x"4b",x"71",x"0e",x"5c"),
   827 => (x"f0",x"fe",x"4c",x"c0"),
   828 => (x"99",x"49",x"70",x"87"),
   829 => (x"87",x"f9",x"c0",x"02"),
   830 => (x"02",x"a9",x"ec",x"c0"),
   831 => (x"c0",x"87",x"f2",x"c0"),
   832 => (x"c0",x"02",x"a9",x"fb"),
   833 => (x"66",x"cc",x"87",x"eb"),
   834 => (x"c7",x"03",x"ac",x"b7"),
   835 => (x"02",x"66",x"d0",x"87"),
   836 => (x"53",x"71",x"87",x"c2"),
   837 => (x"c2",x"02",x"99",x"71"),
   838 => (x"fe",x"84",x"c1",x"87"),
   839 => (x"49",x"70",x"87",x"c3"),
   840 => (x"87",x"cd",x"02",x"99"),
   841 => (x"02",x"a9",x"ec",x"c0"),
   842 => (x"fb",x"c0",x"87",x"c7"),
   843 => (x"d5",x"ff",x"05",x"a9"),
   844 => (x"02",x"66",x"d0",x"87"),
   845 => (x"97",x"c0",x"87",x"c3"),
   846 => (x"a9",x"ec",x"c0",x"7b"),
   847 => (x"74",x"87",x"c4",x"05"),
   848 => (x"74",x"87",x"c5",x"4a"),
   849 => (x"8a",x"0a",x"c0",x"4a"),
   850 => (x"87",x"c2",x"48",x"72"),
   851 => (x"4c",x"26",x"4d",x"26"),
   852 => (x"4f",x"26",x"4b",x"26"),
   853 => (x"87",x"c9",x"fd",x"1e"),
   854 => (x"f0",x"c0",x"49",x"70"),
   855 => (x"ca",x"04",x"a9",x"b7"),
   856 => (x"b7",x"f9",x"c0",x"87"),
   857 => (x"87",x"c3",x"01",x"a9"),
   858 => (x"c1",x"89",x"f0",x"c0"),
   859 => (x"04",x"a9",x"b7",x"c1"),
   860 => (x"da",x"c1",x"87",x"ca"),
   861 => (x"c3",x"01",x"a9",x"b7"),
   862 => (x"89",x"f7",x"c0",x"87"),
   863 => (x"4f",x"26",x"48",x"71"),
   864 => (x"5c",x"5b",x"5e",x"0e"),
   865 => (x"ff",x"4a",x"71",x"0e"),
   866 => (x"49",x"72",x"4c",x"d4"),
   867 => (x"70",x"87",x"ea",x"c0"),
   868 => (x"c2",x"02",x"9b",x"4b"),
   869 => (x"ff",x"8b",x"c1",x"87"),
   870 => (x"c5",x"c8",x"48",x"d0"),
   871 => (x"7c",x"d5",x"c1",x"78"),
   872 => (x"31",x"c6",x"49",x"73"),
   873 => (x"97",x"c3",x"e3",x"c2"),
   874 => (x"71",x"48",x"4a",x"bf"),
   875 => (x"ff",x"7c",x"70",x"b0"),
   876 => (x"78",x"c4",x"48",x"d0"),
   877 => (x"d5",x"fe",x"48",x"73"),
   878 => (x"5b",x"5e",x"0e",x"87"),
   879 => (x"f8",x"0e",x"5d",x"5c"),
   880 => (x"c0",x"4b",x"71",x"86"),
   881 => (x"e0",x"fa",x"c0",x"7e"),
   882 => (x"df",x"49",x"bf",x"97"),
   883 => (x"ee",x"c0",x"05",x"a9"),
   884 => (x"49",x"a3",x"c8",x"87"),
   885 => (x"c1",x"49",x"69",x"97"),
   886 => (x"dd",x"05",x"a9",x"c3"),
   887 => (x"49",x"a3",x"c9",x"87"),
   888 => (x"c1",x"49",x"69",x"97"),
   889 => (x"d1",x"05",x"a9",x"c6"),
   890 => (x"49",x"a3",x"ca",x"87"),
   891 => (x"c1",x"49",x"69",x"97"),
   892 => (x"c5",x"05",x"a9",x"c7"),
   893 => (x"c2",x"48",x"c1",x"87"),
   894 => (x"48",x"c0",x"87",x"e1"),
   895 => (x"fa",x"87",x"dc",x"c2"),
   896 => (x"4c",x"c0",x"87",x"ea"),
   897 => (x"97",x"e0",x"fa",x"c0"),
   898 => (x"a9",x"c0",x"49",x"bf"),
   899 => (x"fa",x"87",x"cf",x"04"),
   900 => (x"84",x"c1",x"87",x"ff"),
   901 => (x"97",x"e0",x"fa",x"c0"),
   902 => (x"06",x"ac",x"49",x"bf"),
   903 => (x"fa",x"c0",x"87",x"f1"),
   904 => (x"02",x"bf",x"97",x"e0"),
   905 => (x"f8",x"f9",x"87",x"cf"),
   906 => (x"99",x"49",x"70",x"87"),
   907 => (x"c0",x"87",x"c6",x"02"),
   908 => (x"f1",x"05",x"a9",x"ec"),
   909 => (x"f9",x"4c",x"c0",x"87"),
   910 => (x"4d",x"70",x"87",x"e7"),
   911 => (x"c8",x"87",x"e2",x"f9"),
   912 => (x"dc",x"f9",x"58",x"a6"),
   913 => (x"c1",x"4a",x"70",x"87"),
   914 => (x"49",x"a3",x"c8",x"84"),
   915 => (x"ad",x"49",x"69",x"97"),
   916 => (x"c0",x"87",x"c7",x"02"),
   917 => (x"c0",x"05",x"ad",x"ff"),
   918 => (x"a3",x"c9",x"87",x"e7"),
   919 => (x"49",x"69",x"97",x"49"),
   920 => (x"02",x"a9",x"66",x"c4"),
   921 => (x"c0",x"48",x"87",x"c7"),
   922 => (x"d4",x"05",x"a8",x"ff"),
   923 => (x"49",x"a3",x"ca",x"87"),
   924 => (x"aa",x"49",x"69",x"97"),
   925 => (x"c0",x"87",x"c6",x"02"),
   926 => (x"c4",x"05",x"aa",x"ff"),
   927 => (x"d0",x"7e",x"c1",x"87"),
   928 => (x"ad",x"ec",x"c0",x"87"),
   929 => (x"c0",x"87",x"c6",x"02"),
   930 => (x"c4",x"05",x"ad",x"fb"),
   931 => (x"c1",x"4c",x"c0",x"87"),
   932 => (x"fe",x"02",x"6e",x"7e"),
   933 => (x"ef",x"f8",x"87",x"e1"),
   934 => (x"f8",x"48",x"74",x"87"),
   935 => (x"87",x"ec",x"fa",x"8e"),
   936 => (x"5b",x"5e",x"0e",x"00"),
   937 => (x"1e",x"0e",x"5d",x"5c"),
   938 => (x"4c",x"c0",x"4b",x"71"),
   939 => (x"c0",x"04",x"ab",x"4d"),
   940 => (x"f6",x"c0",x"87",x"e8"),
   941 => (x"9d",x"75",x"1e",x"f9"),
   942 => (x"c0",x"87",x"c4",x"02"),
   943 => (x"c1",x"87",x"c2",x"4a"),
   944 => (x"ef",x"49",x"72",x"4a"),
   945 => (x"86",x"c4",x"87",x"e6"),
   946 => (x"84",x"c1",x"7e",x"70"),
   947 => (x"87",x"c2",x"05",x"6e"),
   948 => (x"85",x"c1",x"4c",x"73"),
   949 => (x"ff",x"06",x"ac",x"73"),
   950 => (x"48",x"6e",x"87",x"d8"),
   951 => (x"26",x"4d",x"26",x"26"),
   952 => (x"26",x"4b",x"26",x"4c"),
   953 => (x"5b",x"5e",x"0e",x"4f"),
   954 => (x"1e",x"0e",x"5d",x"5c"),
   955 => (x"de",x"49",x"4c",x"71"),
   956 => (x"fd",x"f3",x"c2",x"91"),
   957 => (x"97",x"85",x"71",x"4d"),
   958 => (x"dd",x"c1",x"02",x"6d"),
   959 => (x"e8",x"f3",x"c2",x"87"),
   960 => (x"82",x"74",x"4a",x"bf"),
   961 => (x"d8",x"fe",x"49",x"72"),
   962 => (x"6e",x"7e",x"70",x"87"),
   963 => (x"87",x"f3",x"c0",x"02"),
   964 => (x"4b",x"f0",x"f3",x"c2"),
   965 => (x"49",x"cb",x"4a",x"6e"),
   966 => (x"87",x"cc",x"c6",x"ff"),
   967 => (x"93",x"cb",x"4b",x"74"),
   968 => (x"83",x"d9",x"e2",x"c1"),
   969 => (x"fd",x"c0",x"83",x"c4"),
   970 => (x"49",x"74",x"7b",x"de"),
   971 => (x"87",x"d0",x"c7",x"c1"),
   972 => (x"f3",x"c2",x"7b",x"75"),
   973 => (x"49",x"bf",x"97",x"fc"),
   974 => (x"f0",x"f3",x"c2",x"1e"),
   975 => (x"e6",x"e4",x"c1",x"49"),
   976 => (x"74",x"86",x"c4",x"87"),
   977 => (x"f7",x"c6",x"c1",x"49"),
   978 => (x"c1",x"49",x"c0",x"87"),
   979 => (x"c2",x"87",x"d6",x"c8"),
   980 => (x"c0",x"48",x"e4",x"f3"),
   981 => (x"df",x"49",x"c1",x"78"),
   982 => (x"fd",x"26",x"87",x"fd"),
   983 => (x"6f",x"4c",x"87",x"ff"),
   984 => (x"6e",x"69",x"64",x"61"),
   985 => (x"2e",x"2e",x"2e",x"67"),
   986 => (x"5b",x"5e",x"0e",x"00"),
   987 => (x"4b",x"71",x"0e",x"5c"),
   988 => (x"e8",x"f3",x"c2",x"4a"),
   989 => (x"49",x"72",x"82",x"bf"),
   990 => (x"70",x"87",x"e6",x"fc"),
   991 => (x"c4",x"02",x"9c",x"4c"),
   992 => (x"ef",x"eb",x"49",x"87"),
   993 => (x"e8",x"f3",x"c2",x"87"),
   994 => (x"c1",x"78",x"c0",x"48"),
   995 => (x"87",x"c7",x"df",x"49"),
   996 => (x"0e",x"87",x"cc",x"fd"),
   997 => (x"5d",x"5c",x"5b",x"5e"),
   998 => (x"c2",x"86",x"f4",x"0e"),
   999 => (x"c0",x"4d",x"f2",x"e6"),
  1000 => (x"48",x"a6",x"c4",x"4c"),
  1001 => (x"f3",x"c2",x"78",x"c0"),
  1002 => (x"c0",x"49",x"bf",x"e8"),
  1003 => (x"c1",x"c1",x"06",x"a9"),
  1004 => (x"f2",x"e6",x"c2",x"87"),
  1005 => (x"c0",x"02",x"98",x"48"),
  1006 => (x"f6",x"c0",x"87",x"f8"),
  1007 => (x"66",x"c8",x"1e",x"f9"),
  1008 => (x"c4",x"87",x"c7",x"02"),
  1009 => (x"78",x"c0",x"48",x"a6"),
  1010 => (x"a6",x"c4",x"87",x"c5"),
  1011 => (x"c4",x"78",x"c1",x"48"),
  1012 => (x"d7",x"eb",x"49",x"66"),
  1013 => (x"70",x"86",x"c4",x"87"),
  1014 => (x"c4",x"84",x"c1",x"4d"),
  1015 => (x"80",x"c1",x"48",x"66"),
  1016 => (x"c2",x"58",x"a6",x"c8"),
  1017 => (x"49",x"bf",x"e8",x"f3"),
  1018 => (x"87",x"c6",x"03",x"ac"),
  1019 => (x"ff",x"05",x"9d",x"75"),
  1020 => (x"4c",x"c0",x"87",x"c8"),
  1021 => (x"c3",x"02",x"9d",x"75"),
  1022 => (x"f6",x"c0",x"87",x"e0"),
  1023 => (x"66",x"c8",x"1e",x"f9"),
  1024 => (x"cc",x"87",x"c7",x"02"),
  1025 => (x"78",x"c0",x"48",x"a6"),
  1026 => (x"a6",x"cc",x"87",x"c5"),
  1027 => (x"cc",x"78",x"c1",x"48"),
  1028 => (x"d7",x"ea",x"49",x"66"),
  1029 => (x"70",x"86",x"c4",x"87"),
  1030 => (x"c2",x"02",x"6e",x"7e"),
  1031 => (x"49",x"6e",x"87",x"e9"),
  1032 => (x"69",x"97",x"81",x"cb"),
  1033 => (x"02",x"99",x"d0",x"49"),
  1034 => (x"c0",x"87",x"d6",x"c1"),
  1035 => (x"74",x"4a",x"e9",x"fd"),
  1036 => (x"c1",x"91",x"cb",x"49"),
  1037 => (x"72",x"81",x"d9",x"e2"),
  1038 => (x"c3",x"81",x"c8",x"79"),
  1039 => (x"49",x"74",x"51",x"ff"),
  1040 => (x"f3",x"c2",x"91",x"de"),
  1041 => (x"85",x"71",x"4d",x"fd"),
  1042 => (x"7d",x"97",x"c1",x"c2"),
  1043 => (x"c0",x"49",x"a5",x"c1"),
  1044 => (x"ef",x"c2",x"51",x"e0"),
  1045 => (x"02",x"bf",x"97",x"c2"),
  1046 => (x"84",x"c1",x"87",x"d2"),
  1047 => (x"c2",x"4b",x"a5",x"c2"),
  1048 => (x"db",x"4a",x"c2",x"ef"),
  1049 => (x"ff",x"c0",x"ff",x"49"),
  1050 => (x"87",x"db",x"c1",x"87"),
  1051 => (x"c0",x"49",x"a5",x"cd"),
  1052 => (x"c2",x"84",x"c1",x"51"),
  1053 => (x"4a",x"6e",x"4b",x"a5"),
  1054 => (x"c0",x"ff",x"49",x"cb"),
  1055 => (x"c6",x"c1",x"87",x"ea"),
  1056 => (x"e5",x"fb",x"c0",x"87"),
  1057 => (x"cb",x"49",x"74",x"4a"),
  1058 => (x"d9",x"e2",x"c1",x"91"),
  1059 => (x"c2",x"79",x"72",x"81"),
  1060 => (x"bf",x"97",x"c2",x"ef"),
  1061 => (x"74",x"87",x"d8",x"02"),
  1062 => (x"c1",x"91",x"de",x"49"),
  1063 => (x"fd",x"f3",x"c2",x"84"),
  1064 => (x"c2",x"83",x"71",x"4b"),
  1065 => (x"dd",x"4a",x"c2",x"ef"),
  1066 => (x"fb",x"ff",x"fe",x"49"),
  1067 => (x"74",x"87",x"d8",x"87"),
  1068 => (x"c2",x"93",x"de",x"4b"),
  1069 => (x"cb",x"83",x"fd",x"f3"),
  1070 => (x"51",x"c0",x"49",x"a3"),
  1071 => (x"6e",x"73",x"84",x"c1"),
  1072 => (x"fe",x"49",x"cb",x"4a"),
  1073 => (x"c4",x"87",x"e1",x"ff"),
  1074 => (x"80",x"c1",x"48",x"66"),
  1075 => (x"c7",x"58",x"a6",x"c8"),
  1076 => (x"c5",x"c0",x"03",x"ac"),
  1077 => (x"fc",x"05",x"6e",x"87"),
  1078 => (x"48",x"74",x"87",x"e0"),
  1079 => (x"fc",x"f7",x"8e",x"f4"),
  1080 => (x"1e",x"73",x"1e",x"87"),
  1081 => (x"cb",x"49",x"4b",x"71"),
  1082 => (x"d9",x"e2",x"c1",x"91"),
  1083 => (x"4a",x"a1",x"c8",x"81"),
  1084 => (x"48",x"c3",x"e3",x"c2"),
  1085 => (x"a1",x"c9",x"50",x"12"),
  1086 => (x"e0",x"fa",x"c0",x"4a"),
  1087 => (x"ca",x"50",x"12",x"48"),
  1088 => (x"fc",x"f3",x"c2",x"81"),
  1089 => (x"c2",x"50",x"11",x"48"),
  1090 => (x"bf",x"97",x"fc",x"f3"),
  1091 => (x"49",x"c0",x"1e",x"49"),
  1092 => (x"87",x"d3",x"dd",x"c1"),
  1093 => (x"48",x"e4",x"f3",x"c2"),
  1094 => (x"49",x"c1",x"78",x"de"),
  1095 => (x"26",x"87",x"f8",x"d8"),
  1096 => (x"1e",x"87",x"fe",x"f6"),
  1097 => (x"cb",x"49",x"4a",x"71"),
  1098 => (x"d9",x"e2",x"c1",x"91"),
  1099 => (x"11",x"81",x"c8",x"81"),
  1100 => (x"e8",x"f3",x"c2",x"48"),
  1101 => (x"e8",x"f3",x"c2",x"58"),
  1102 => (x"c1",x"78",x"c0",x"48"),
  1103 => (x"87",x"d7",x"d8",x"49"),
  1104 => (x"c0",x"1e",x"4f",x"26"),
  1105 => (x"dc",x"c0",x"c1",x"49"),
  1106 => (x"1e",x"4f",x"26",x"87"),
  1107 => (x"d2",x"02",x"99",x"71"),
  1108 => (x"ee",x"e3",x"c1",x"87"),
  1109 => (x"f7",x"50",x"c0",x"48"),
  1110 => (x"e3",x"c4",x"c1",x"80"),
  1111 => (x"c7",x"e2",x"c1",x"40"),
  1112 => (x"c1",x"87",x"ce",x"78"),
  1113 => (x"c1",x"48",x"ea",x"e3"),
  1114 => (x"fc",x"78",x"e8",x"e1"),
  1115 => (x"c2",x"c5",x"c1",x"80"),
  1116 => (x"0e",x"4f",x"26",x"78"),
  1117 => (x"0e",x"5c",x"5b",x"5e"),
  1118 => (x"cb",x"4a",x"4c",x"71"),
  1119 => (x"d9",x"e2",x"c1",x"92"),
  1120 => (x"49",x"a2",x"c8",x"82"),
  1121 => (x"97",x"4b",x"a2",x"c9"),
  1122 => (x"97",x"1e",x"4b",x"6b"),
  1123 => (x"ca",x"1e",x"49",x"69"),
  1124 => (x"c0",x"49",x"12",x"82"),
  1125 => (x"c0",x"87",x"d7",x"eb"),
  1126 => (x"87",x"fb",x"d6",x"49"),
  1127 => (x"fd",x"c0",x"49",x"74"),
  1128 => (x"8e",x"f8",x"87",x"de"),
  1129 => (x"1e",x"87",x"f8",x"f4"),
  1130 => (x"4b",x"71",x"1e",x"73"),
  1131 => (x"87",x"c3",x"ff",x"49"),
  1132 => (x"fe",x"fe",x"49",x"73"),
  1133 => (x"87",x"e9",x"f4",x"87"),
  1134 => (x"71",x"1e",x"73",x"1e"),
  1135 => (x"4a",x"a3",x"c6",x"4b"),
  1136 => (x"c1",x"87",x"dc",x"02"),
  1137 => (x"e4",x"c0",x"02",x"8a"),
  1138 => (x"c1",x"02",x"8a",x"87"),
  1139 => (x"02",x"8a",x"87",x"e8"),
  1140 => (x"8a",x"87",x"ca",x"c1"),
  1141 => (x"87",x"ef",x"c0",x"02"),
  1142 => (x"87",x"d9",x"02",x"8a"),
  1143 => (x"c2",x"87",x"e9",x"c1"),
  1144 => (x"df",x"48",x"e4",x"f3"),
  1145 => (x"d5",x"49",x"c1",x"78"),
  1146 => (x"e6",x"c1",x"87",x"ed"),
  1147 => (x"fc",x"49",x"c7",x"87"),
  1148 => (x"de",x"c1",x"87",x"f1"),
  1149 => (x"e8",x"f3",x"c2",x"87"),
  1150 => (x"cb",x"c1",x"02",x"bf"),
  1151 => (x"88",x"c1",x"48",x"87"),
  1152 => (x"58",x"ec",x"f3",x"c2"),
  1153 => (x"c2",x"87",x"c1",x"c1"),
  1154 => (x"02",x"bf",x"ec",x"f3"),
  1155 => (x"c2",x"87",x"f9",x"c0"),
  1156 => (x"48",x"bf",x"e8",x"f3"),
  1157 => (x"f3",x"c2",x"80",x"c1"),
  1158 => (x"eb",x"c0",x"58",x"ec"),
  1159 => (x"e8",x"f3",x"c2",x"87"),
  1160 => (x"89",x"c6",x"49",x"bf"),
  1161 => (x"59",x"ec",x"f3",x"c2"),
  1162 => (x"03",x"a9",x"b7",x"c0"),
  1163 => (x"f3",x"c2",x"87",x"da"),
  1164 => (x"78",x"c0",x"48",x"e8"),
  1165 => (x"f3",x"c2",x"87",x"d2"),
  1166 => (x"cb",x"02",x"bf",x"ec"),
  1167 => (x"e8",x"f3",x"c2",x"87"),
  1168 => (x"80",x"c6",x"48",x"bf"),
  1169 => (x"58",x"ec",x"f3",x"c2"),
  1170 => (x"ca",x"d4",x"49",x"c0"),
  1171 => (x"c0",x"49",x"73",x"87"),
  1172 => (x"f2",x"87",x"ed",x"fa"),
  1173 => (x"5e",x"0e",x"87",x"cb"),
  1174 => (x"71",x"0e",x"5c",x"5b"),
  1175 => (x"1e",x"66",x"cc",x"4c"),
  1176 => (x"93",x"cb",x"4b",x"74"),
  1177 => (x"83",x"d9",x"e2",x"c1"),
  1178 => (x"6a",x"4a",x"a3",x"c4"),
  1179 => (x"c7",x"f9",x"fe",x"49"),
  1180 => (x"e1",x"c3",x"c1",x"87"),
  1181 => (x"49",x"a3",x"c8",x"7b"),
  1182 => (x"c9",x"51",x"66",x"d4"),
  1183 => (x"66",x"d8",x"49",x"a3"),
  1184 => (x"49",x"a3",x"ca",x"51"),
  1185 => (x"26",x"51",x"66",x"dc"),
  1186 => (x"0e",x"87",x"d4",x"f1"),
  1187 => (x"5d",x"5c",x"5b",x"5e"),
  1188 => (x"86",x"d0",x"ff",x"0e"),
  1189 => (x"c8",x"59",x"a6",x"d8"),
  1190 => (x"78",x"c0",x"48",x"a6"),
  1191 => (x"c4",x"c1",x"80",x"fc"),
  1192 => (x"80",x"c8",x"78",x"66"),
  1193 => (x"80",x"c4",x"78",x"c1"),
  1194 => (x"f3",x"c2",x"78",x"c1"),
  1195 => (x"78",x"c1",x"48",x"ec"),
  1196 => (x"bf",x"e4",x"f3",x"c2"),
  1197 => (x"de",x"48",x"6e",x"7e"),
  1198 => (x"87",x"cb",x"05",x"a8"),
  1199 => (x"70",x"87",x"d4",x"f3"),
  1200 => (x"59",x"a6",x"cc",x"49"),
  1201 => (x"6e",x"87",x"f8",x"d0"),
  1202 => (x"05",x"a8",x"df",x"48"),
  1203 => (x"c1",x"87",x"ee",x"c1"),
  1204 => (x"c4",x"49",x"66",x"c0"),
  1205 => (x"c1",x"7e",x"69",x"81"),
  1206 => (x"6e",x"48",x"f4",x"dc"),
  1207 => (x"4a",x"a1",x"d0",x"49"),
  1208 => (x"aa",x"71",x"41",x"20"),
  1209 => (x"c1",x"87",x"f9",x"05"),
  1210 => (x"c1",x"4a",x"e1",x"c3"),
  1211 => (x"7a",x"0a",x"66",x"c0"),
  1212 => (x"66",x"c0",x"c1",x"0a"),
  1213 => (x"df",x"81",x"c9",x"49"),
  1214 => (x"66",x"c0",x"c1",x"51"),
  1215 => (x"c1",x"81",x"ca",x"49"),
  1216 => (x"c0",x"c1",x"51",x"d3"),
  1217 => (x"81",x"cb",x"49",x"66"),
  1218 => (x"c4",x"4b",x"a1",x"c4"),
  1219 => (x"78",x"6b",x"48",x"a6"),
  1220 => (x"1e",x"72",x"1e",x"71"),
  1221 => (x"48",x"c4",x"dd",x"c1"),
  1222 => (x"d0",x"49",x"66",x"cc"),
  1223 => (x"41",x"20",x"4a",x"a1"),
  1224 => (x"f9",x"05",x"aa",x"71"),
  1225 => (x"26",x"4a",x"26",x"87"),
  1226 => (x"c9",x"79",x"72",x"49"),
  1227 => (x"52",x"df",x"4a",x"a1"),
  1228 => (x"d4",x"c1",x"81",x"ca"),
  1229 => (x"48",x"a6",x"c8",x"51"),
  1230 => (x"c2",x"cf",x"78",x"c2"),
  1231 => (x"87",x"ec",x"e5",x"87"),
  1232 => (x"e5",x"87",x"ce",x"e6"),
  1233 => (x"4c",x"70",x"87",x"db"),
  1234 => (x"02",x"ac",x"fb",x"c0"),
  1235 => (x"d4",x"87",x"d0",x"c1"),
  1236 => (x"c2",x"c1",x"05",x"66"),
  1237 => (x"1e",x"1e",x"c0",x"87"),
  1238 => (x"e4",x"c1",x"1e",x"c1"),
  1239 => (x"49",x"c0",x"1e",x"cc"),
  1240 => (x"c1",x"87",x"f3",x"fb"),
  1241 => (x"c4",x"4a",x"66",x"d0"),
  1242 => (x"c7",x"49",x"6a",x"82"),
  1243 => (x"c1",x"51",x"74",x"81"),
  1244 => (x"6a",x"1e",x"d8",x"1e"),
  1245 => (x"e5",x"81",x"c8",x"49"),
  1246 => (x"86",x"d8",x"87",x"eb"),
  1247 => (x"48",x"66",x"c4",x"c1"),
  1248 => (x"c7",x"01",x"a8",x"c0"),
  1249 => (x"48",x"a6",x"c8",x"87"),
  1250 => (x"87",x"ce",x"78",x"c1"),
  1251 => (x"48",x"66",x"c4",x"c1"),
  1252 => (x"a6",x"c8",x"88",x"c1"),
  1253 => (x"e4",x"87",x"c3",x"58"),
  1254 => (x"a6",x"cc",x"87",x"f7"),
  1255 => (x"74",x"78",x"c2",x"48"),
  1256 => (x"d6",x"cd",x"02",x"9c"),
  1257 => (x"48",x"66",x"c8",x"87"),
  1258 => (x"a8",x"66",x"c8",x"c1"),
  1259 => (x"87",x"cb",x"cd",x"03"),
  1260 => (x"c0",x"48",x"a6",x"d8"),
  1261 => (x"87",x"e9",x"e3",x"78"),
  1262 => (x"d0",x"c1",x"4c",x"70"),
  1263 => (x"d6",x"c2",x"05",x"ac"),
  1264 => (x"7e",x"66",x"d8",x"87"),
  1265 => (x"70",x"87",x"cd",x"e6"),
  1266 => (x"59",x"a6",x"dc",x"49"),
  1267 => (x"70",x"87",x"d2",x"e3"),
  1268 => (x"ac",x"ec",x"c0",x"4c"),
  1269 => (x"87",x"ea",x"c1",x"05"),
  1270 => (x"cb",x"49",x"66",x"c8"),
  1271 => (x"66",x"c0",x"c1",x"91"),
  1272 => (x"4a",x"a1",x"c4",x"81"),
  1273 => (x"a1",x"c8",x"4d",x"6a"),
  1274 => (x"52",x"66",x"d8",x"4a"),
  1275 => (x"79",x"e3",x"c4",x"c1"),
  1276 => (x"70",x"87",x"ee",x"e2"),
  1277 => (x"d8",x"02",x"9c",x"4c"),
  1278 => (x"ac",x"fb",x"c0",x"87"),
  1279 => (x"74",x"87",x"d2",x"02"),
  1280 => (x"87",x"dd",x"e2",x"55"),
  1281 => (x"02",x"9c",x"4c",x"70"),
  1282 => (x"fb",x"c0",x"87",x"c7"),
  1283 => (x"ee",x"ff",x"05",x"ac"),
  1284 => (x"55",x"e0",x"c0",x"87"),
  1285 => (x"c0",x"55",x"c1",x"c2"),
  1286 => (x"66",x"d4",x"7d",x"97"),
  1287 => (x"05",x"a9",x"6e",x"49"),
  1288 => (x"66",x"c8",x"87",x"db"),
  1289 => (x"a8",x"66",x"c4",x"48"),
  1290 => (x"c8",x"87",x"ca",x"04"),
  1291 => (x"80",x"c1",x"48",x"66"),
  1292 => (x"c8",x"58",x"a6",x"cc"),
  1293 => (x"48",x"66",x"c4",x"87"),
  1294 => (x"a6",x"c8",x"88",x"c1"),
  1295 => (x"87",x"e1",x"e1",x"58"),
  1296 => (x"d0",x"c1",x"4c",x"70"),
  1297 => (x"87",x"c8",x"05",x"ac"),
  1298 => (x"c1",x"48",x"66",x"d0"),
  1299 => (x"58",x"a6",x"d4",x"80"),
  1300 => (x"02",x"ac",x"d0",x"c1"),
  1301 => (x"dc",x"87",x"ea",x"fd"),
  1302 => (x"66",x"d4",x"48",x"a6"),
  1303 => (x"48",x"66",x"d8",x"78"),
  1304 => (x"05",x"a8",x"66",x"dc"),
  1305 => (x"c0",x"87",x"e6",x"c9"),
  1306 => (x"c0",x"48",x"a6",x"e0"),
  1307 => (x"80",x"c4",x"78",x"f0"),
  1308 => (x"c4",x"78",x"66",x"cc"),
  1309 => (x"7e",x"78",x"c0",x"80"),
  1310 => (x"fb",x"c0",x"48",x"74"),
  1311 => (x"a6",x"f0",x"c0",x"88"),
  1312 => (x"02",x"98",x"70",x"58"),
  1313 => (x"48",x"87",x"e1",x"c8"),
  1314 => (x"f0",x"c0",x"88",x"cb"),
  1315 => (x"98",x"70",x"58",x"a6"),
  1316 => (x"87",x"e9",x"c0",x"02"),
  1317 => (x"c0",x"88",x"c9",x"48"),
  1318 => (x"70",x"58",x"a6",x"f0"),
  1319 => (x"e9",x"c3",x"02",x"98"),
  1320 => (x"88",x"c4",x"48",x"87"),
  1321 => (x"58",x"a6",x"f0",x"c0"),
  1322 => (x"de",x"02",x"98",x"70"),
  1323 => (x"88",x"c1",x"48",x"87"),
  1324 => (x"58",x"a6",x"f0",x"c0"),
  1325 => (x"c3",x"02",x"98",x"70"),
  1326 => (x"e5",x"c7",x"87",x"d0"),
  1327 => (x"a6",x"e0",x"c0",x"87"),
  1328 => (x"cc",x"78",x"c0",x"48"),
  1329 => (x"80",x"c1",x"48",x"66"),
  1330 => (x"ff",x"58",x"a6",x"d0"),
  1331 => (x"70",x"87",x"d2",x"df"),
  1332 => (x"ac",x"ec",x"c0",x"4c"),
  1333 => (x"c0",x"87",x"d7",x"02"),
  1334 => (x"c0",x"02",x"66",x"e0"),
  1335 => (x"e4",x"c0",x"87",x"c7"),
  1336 => (x"c9",x"c0",x"5c",x"a6"),
  1337 => (x"c0",x"48",x"74",x"87"),
  1338 => (x"e8",x"c0",x"88",x"f0"),
  1339 => (x"ec",x"c0",x"58",x"a6"),
  1340 => (x"cd",x"c0",x"02",x"ac"),
  1341 => (x"e8",x"de",x"ff",x"87"),
  1342 => (x"c0",x"4c",x"70",x"87"),
  1343 => (x"ff",x"05",x"ac",x"ec"),
  1344 => (x"e0",x"c0",x"87",x"f3"),
  1345 => (x"66",x"d4",x"1e",x"66"),
  1346 => (x"ec",x"c0",x"1e",x"49"),
  1347 => (x"e4",x"c1",x"1e",x"66"),
  1348 => (x"66",x"d8",x"1e",x"cc"),
  1349 => (x"87",x"fe",x"f4",x"49"),
  1350 => (x"1e",x"ca",x"1e",x"c0"),
  1351 => (x"49",x"66",x"e0",x"c0"),
  1352 => (x"d8",x"c1",x"91",x"cb"),
  1353 => (x"a6",x"d8",x"81",x"66"),
  1354 => (x"78",x"a1",x"c4",x"48"),
  1355 => (x"49",x"bf",x"66",x"d8"),
  1356 => (x"87",x"f1",x"de",x"ff"),
  1357 => (x"b7",x"c0",x"86",x"d8"),
  1358 => (x"c8",x"c1",x"06",x"a8"),
  1359 => (x"de",x"1e",x"c1",x"87"),
  1360 => (x"bf",x"66",x"c8",x"1e"),
  1361 => (x"dc",x"de",x"ff",x"49"),
  1362 => (x"70",x"86",x"c8",x"87"),
  1363 => (x"08",x"c0",x"48",x"49"),
  1364 => (x"a6",x"e4",x"c0",x"88"),
  1365 => (x"a8",x"b7",x"c0",x"58"),
  1366 => (x"87",x"e9",x"c0",x"06"),
  1367 => (x"48",x"66",x"e0",x"c0"),
  1368 => (x"03",x"a8",x"b7",x"dd"),
  1369 => (x"bf",x"6e",x"87",x"df"),
  1370 => (x"66",x"e0",x"c0",x"49"),
  1371 => (x"51",x"e0",x"c0",x"81"),
  1372 => (x"81",x"c1",x"49",x"66"),
  1373 => (x"c2",x"81",x"bf",x"6e"),
  1374 => (x"e0",x"c0",x"51",x"c1"),
  1375 => (x"81",x"c2",x"49",x"66"),
  1376 => (x"c0",x"81",x"bf",x"6e"),
  1377 => (x"c4",x"7e",x"c1",x"51"),
  1378 => (x"df",x"ff",x"87",x"de"),
  1379 => (x"e4",x"c0",x"87",x"c6"),
  1380 => (x"de",x"ff",x"58",x"a6"),
  1381 => (x"e8",x"c0",x"87",x"fe"),
  1382 => (x"ec",x"c0",x"58",x"a6"),
  1383 => (x"cb",x"c0",x"05",x"a8"),
  1384 => (x"a6",x"e4",x"c0",x"87"),
  1385 => (x"66",x"e0",x"c0",x"48"),
  1386 => (x"87",x"c4",x"c0",x"78"),
  1387 => (x"87",x"f1",x"db",x"ff"),
  1388 => (x"cb",x"49",x"66",x"c8"),
  1389 => (x"66",x"c0",x"c1",x"91"),
  1390 => (x"70",x"80",x"71",x"48"),
  1391 => (x"c8",x"4a",x"6e",x"7e"),
  1392 => (x"ca",x"49",x"6e",x"82"),
  1393 => (x"66",x"e0",x"c0",x"81"),
  1394 => (x"66",x"e4",x"c0",x"51"),
  1395 => (x"c0",x"81",x"c1",x"49"),
  1396 => (x"c1",x"89",x"66",x"e0"),
  1397 => (x"70",x"30",x"71",x"48"),
  1398 => (x"71",x"89",x"c1",x"49"),
  1399 => (x"f7",x"c2",x"7a",x"97"),
  1400 => (x"c0",x"49",x"bf",x"d9"),
  1401 => (x"97",x"29",x"66",x"e0"),
  1402 => (x"71",x"48",x"4a",x"6a"),
  1403 => (x"a6",x"f0",x"c0",x"98"),
  1404 => (x"c4",x"49",x"6e",x"58"),
  1405 => (x"dc",x"4d",x"69",x"81"),
  1406 => (x"66",x"d8",x"48",x"66"),
  1407 => (x"c8",x"c0",x"02",x"a8"),
  1408 => (x"48",x"a6",x"d8",x"87"),
  1409 => (x"c5",x"c0",x"78",x"c0"),
  1410 => (x"48",x"a6",x"d8",x"87"),
  1411 => (x"66",x"d8",x"78",x"c1"),
  1412 => (x"1e",x"e0",x"c0",x"1e"),
  1413 => (x"db",x"ff",x"49",x"75"),
  1414 => (x"86",x"c8",x"87",x"cb"),
  1415 => (x"b7",x"c0",x"4c",x"70"),
  1416 => (x"d4",x"c1",x"06",x"ac"),
  1417 => (x"c0",x"85",x"74",x"87"),
  1418 => (x"89",x"74",x"49",x"e0"),
  1419 => (x"dd",x"c1",x"4b",x"75"),
  1420 => (x"fe",x"71",x"4a",x"d4"),
  1421 => (x"c2",x"87",x"f1",x"e9"),
  1422 => (x"66",x"e8",x"c0",x"85"),
  1423 => (x"c0",x"80",x"c1",x"48"),
  1424 => (x"c0",x"58",x"a6",x"ec"),
  1425 => (x"c1",x"49",x"66",x"ec"),
  1426 => (x"02",x"a9",x"70",x"81"),
  1427 => (x"d8",x"87",x"c8",x"c0"),
  1428 => (x"78",x"c0",x"48",x"a6"),
  1429 => (x"d8",x"87",x"c5",x"c0"),
  1430 => (x"78",x"c1",x"48",x"a6"),
  1431 => (x"c2",x"1e",x"66",x"d8"),
  1432 => (x"e0",x"c0",x"49",x"a4"),
  1433 => (x"70",x"88",x"71",x"48"),
  1434 => (x"49",x"75",x"1e",x"49"),
  1435 => (x"87",x"f5",x"d9",x"ff"),
  1436 => (x"b7",x"c0",x"86",x"c8"),
  1437 => (x"c0",x"ff",x"01",x"a8"),
  1438 => (x"66",x"e8",x"c0",x"87"),
  1439 => (x"87",x"d1",x"c0",x"02"),
  1440 => (x"81",x"c9",x"49",x"6e"),
  1441 => (x"51",x"66",x"e8",x"c0"),
  1442 => (x"c5",x"c1",x"48",x"6e"),
  1443 => (x"cc",x"c0",x"78",x"f3"),
  1444 => (x"c9",x"49",x"6e",x"87"),
  1445 => (x"6e",x"51",x"c2",x"81"),
  1446 => (x"e7",x"c6",x"c1",x"48"),
  1447 => (x"c0",x"7e",x"c1",x"78"),
  1448 => (x"d8",x"ff",x"87",x"c6"),
  1449 => (x"4c",x"70",x"87",x"eb"),
  1450 => (x"f5",x"c0",x"02",x"6e"),
  1451 => (x"48",x"66",x"c8",x"87"),
  1452 => (x"04",x"a8",x"66",x"c4"),
  1453 => (x"c8",x"87",x"cb",x"c0"),
  1454 => (x"80",x"c1",x"48",x"66"),
  1455 => (x"c0",x"58",x"a6",x"cc"),
  1456 => (x"66",x"c4",x"87",x"e0"),
  1457 => (x"c8",x"88",x"c1",x"48"),
  1458 => (x"d5",x"c0",x"58",x"a6"),
  1459 => (x"ac",x"c6",x"c1",x"87"),
  1460 => (x"87",x"c8",x"c0",x"05"),
  1461 => (x"c1",x"48",x"66",x"cc"),
  1462 => (x"58",x"a6",x"d0",x"80"),
  1463 => (x"87",x"f1",x"d7",x"ff"),
  1464 => (x"66",x"d0",x"4c",x"70"),
  1465 => (x"d4",x"80",x"c1",x"48"),
  1466 => (x"9c",x"74",x"58",x"a6"),
  1467 => (x"87",x"cb",x"c0",x"02"),
  1468 => (x"c1",x"48",x"66",x"c8"),
  1469 => (x"04",x"a8",x"66",x"c8"),
  1470 => (x"ff",x"87",x"f5",x"f2"),
  1471 => (x"c8",x"87",x"c9",x"d7"),
  1472 => (x"a8",x"c7",x"48",x"66"),
  1473 => (x"87",x"e5",x"c0",x"03"),
  1474 => (x"48",x"ec",x"f3",x"c2"),
  1475 => (x"66",x"c8",x"78",x"c0"),
  1476 => (x"c1",x"91",x"cb",x"49"),
  1477 => (x"c4",x"81",x"66",x"c0"),
  1478 => (x"4a",x"6a",x"4a",x"a1"),
  1479 => (x"c8",x"79",x"52",x"c0"),
  1480 => (x"80",x"c1",x"48",x"66"),
  1481 => (x"c7",x"58",x"a6",x"cc"),
  1482 => (x"db",x"ff",x"04",x"a8"),
  1483 => (x"8e",x"d0",x"ff",x"87"),
  1484 => (x"87",x"e9",x"de",x"ff"),
  1485 => (x"64",x"61",x"6f",x"4c"),
  1486 => (x"74",x"65",x"53",x"20"),
  1487 => (x"67",x"6e",x"69",x"74"),
  1488 => (x"00",x"81",x"20",x"73"),
  1489 => (x"65",x"76",x"61",x"53"),
  1490 => (x"74",x"65",x"53",x"20"),
  1491 => (x"67",x"6e",x"69",x"74"),
  1492 => (x"00",x"81",x"20",x"73"),
  1493 => (x"1e",x"00",x"20",x"3a"),
  1494 => (x"4b",x"71",x"1e",x"73"),
  1495 => (x"87",x"c6",x"02",x"9b"),
  1496 => (x"48",x"e8",x"f3",x"c2"),
  1497 => (x"1e",x"c7",x"78",x"c0"),
  1498 => (x"bf",x"e8",x"f3",x"c2"),
  1499 => (x"e2",x"c1",x"1e",x"49"),
  1500 => (x"f3",x"c2",x"1e",x"d9"),
  1501 => (x"ec",x"49",x"bf",x"e4"),
  1502 => (x"86",x"cc",x"87",x"d1"),
  1503 => (x"bf",x"e4",x"f3",x"c2"),
  1504 => (x"87",x"c7",x"e7",x"49"),
  1505 => (x"c8",x"02",x"9b",x"73"),
  1506 => (x"d9",x"e2",x"c1",x"87"),
  1507 => (x"c1",x"e7",x"c0",x"49"),
  1508 => (x"cc",x"dd",x"ff",x"87"),
  1509 => (x"1e",x"73",x"1e",x"87"),
  1510 => (x"df",x"c1",x"4b",x"c0"),
  1511 => (x"c5",x"c1",x"49",x"c0"),
  1512 => (x"e3",x"c2",x"87",x"fc"),
  1513 => (x"50",x"c0",x"48",x"c3"),
  1514 => (x"bf",x"fc",x"e3",x"c1"),
  1515 => (x"c9",x"ff",x"c0",x"49"),
  1516 => (x"05",x"98",x"70",x"87"),
  1517 => (x"df",x"c1",x"87",x"c4"),
  1518 => (x"48",x"73",x"4b",x"cc"),
  1519 => (x"87",x"e1",x"dc",x"ff"),
  1520 => (x"43",x"49",x"52",x"4f"),
  1521 => (x"20",x"20",x"20",x"20"),
  1522 => (x"00",x"47",x"46",x"43"),
  1523 => (x"20",x"4d",x"4f",x"52"),
  1524 => (x"64",x"61",x"6f",x"6c"),
  1525 => (x"20",x"67",x"6e",x"69"),
  1526 => (x"6c",x"69",x"61",x"66"),
  1527 => (x"1e",x"00",x"64",x"65"),
  1528 => (x"c1",x"87",x"c8",x"c8"),
  1529 => (x"87",x"ef",x"fd",x"49"),
  1530 => (x"87",x"cf",x"eb",x"fe"),
  1531 => (x"cd",x"02",x"98",x"70"),
  1532 => (x"cc",x"f4",x"fe",x"87"),
  1533 => (x"02",x"98",x"70",x"87"),
  1534 => (x"4a",x"c1",x"87",x"c4"),
  1535 => (x"4a",x"c0",x"87",x"c2"),
  1536 => (x"ce",x"05",x"9a",x"72"),
  1537 => (x"c1",x"1e",x"c0",x"87"),
  1538 => (x"c0",x"49",x"ef",x"e0"),
  1539 => (x"c4",x"87",x"f9",x"f3"),
  1540 => (x"c0",x"87",x"fe",x"86"),
  1541 => (x"fa",x"e0",x"c1",x"1e"),
  1542 => (x"eb",x"f3",x"c0",x"49"),
  1543 => (x"fd",x"1e",x"c0",x"87"),
  1544 => (x"49",x"70",x"87",x"f3"),
  1545 => (x"87",x"e0",x"f3",x"c0"),
  1546 => (x"f8",x"87",x"ff",x"c3"),
  1547 => (x"53",x"4f",x"26",x"8e"),
  1548 => (x"61",x"66",x"20",x"44"),
  1549 => (x"64",x"65",x"6c",x"69"),
  1550 => (x"6f",x"42",x"00",x"2e"),
  1551 => (x"6e",x"69",x"74",x"6f"),
  1552 => (x"2e",x"2e",x"2e",x"67"),
  1553 => (x"e8",x"c0",x"1e",x"00"),
  1554 => (x"f7",x"c0",x"87",x"eb"),
  1555 => (x"87",x"f6",x"87",x"c5"),
  1556 => (x"c2",x"1e",x"4f",x"26"),
  1557 => (x"c0",x"48",x"e8",x"f3"),
  1558 => (x"e4",x"f3",x"c2",x"78"),
  1559 => (x"fd",x"78",x"c0",x"48"),
  1560 => (x"87",x"e1",x"87",x"fd"),
  1561 => (x"4f",x"26",x"48",x"c0"),
  1562 => (x"20",x"20",x"20",x"20"),
  1563 => (x"20",x"20",x"20",x"20"),
  1564 => (x"20",x"20",x"20",x"20"),
  1565 => (x"69",x"78",x"45",x"20"),
  1566 => (x"20",x"20",x"20",x"74"),
  1567 => (x"20",x"20",x"20",x"20"),
  1568 => (x"20",x"20",x"20",x"20"),
  1569 => (x"80",x"00",x"81",x"20"),
  1570 => (x"20",x"20",x"20",x"20"),
  1571 => (x"20",x"20",x"20",x"20"),
  1572 => (x"20",x"20",x"20",x"20"),
  1573 => (x"6b",x"63",x"61",x"42"),
  1574 => (x"00",x"11",x"23",x"00"),
  1575 => (x"00",x"2c",x"fd",x"00"),
  1576 => (x"00",x"00",x"00",x"00"),
  1577 => (x"00",x"00",x"11",x"23"),
  1578 => (x"00",x"00",x"2d",x"1b"),
  1579 => (x"23",x"00",x"00",x"00"),
  1580 => (x"39",x"00",x"00",x"11"),
  1581 => (x"00",x"00",x"00",x"2d"),
  1582 => (x"11",x"23",x"00",x"00"),
  1583 => (x"2d",x"57",x"00",x"00"),
  1584 => (x"00",x"00",x"00",x"00"),
  1585 => (x"00",x"11",x"23",x"00"),
  1586 => (x"00",x"2d",x"75",x"00"),
  1587 => (x"00",x"00",x"00",x"00"),
  1588 => (x"00",x"00",x"11",x"23"),
  1589 => (x"00",x"00",x"2d",x"93"),
  1590 => (x"23",x"00",x"00",x"00"),
  1591 => (x"b1",x"00",x"00",x"11"),
  1592 => (x"00",x"00",x"00",x"2d"),
  1593 => (x"11",x"23",x"00",x"00"),
  1594 => (x"00",x"00",x"00",x"00"),
  1595 => (x"00",x"00",x"00",x"00"),
  1596 => (x"00",x"11",x"b8",x"00"),
  1597 => (x"00",x"00",x"00",x"00"),
  1598 => (x"00",x"00",x"00",x"00"),
  1599 => (x"00",x"00",x"19",x"00"),
  1600 => (x"43",x"49",x"52",x"4f"),
  1601 => (x"20",x"20",x"20",x"20"),
  1602 => (x"00",x"4d",x"4f",x"52"),
  1603 => (x"64",x"61",x"6f",x"4c"),
  1604 => (x"00",x"2e",x"2a",x"20"),
  1605 => (x"48",x"f0",x"fe",x"1e"),
  1606 => (x"09",x"cd",x"78",x"c0"),
  1607 => (x"4f",x"26",x"09",x"79"),
  1608 => (x"f0",x"fe",x"1e",x"1e"),
  1609 => (x"26",x"48",x"7e",x"bf"),
  1610 => (x"fe",x"1e",x"4f",x"26"),
  1611 => (x"78",x"c1",x"48",x"f0"),
  1612 => (x"fe",x"1e",x"4f",x"26"),
  1613 => (x"78",x"c0",x"48",x"f0"),
  1614 => (x"71",x"1e",x"4f",x"26"),
  1615 => (x"52",x"52",x"c0",x"4a"),
  1616 => (x"5e",x"0e",x"4f",x"26"),
  1617 => (x"0e",x"5d",x"5c",x"5b"),
  1618 => (x"4d",x"71",x"86",x"f4"),
  1619 => (x"c1",x"7e",x"6d",x"97"),
  1620 => (x"6c",x"97",x"4c",x"a5"),
  1621 => (x"58",x"a6",x"c8",x"48"),
  1622 => (x"66",x"c4",x"48",x"6e"),
  1623 => (x"87",x"c5",x"05",x"a8"),
  1624 => (x"e6",x"c0",x"48",x"ff"),
  1625 => (x"87",x"ca",x"ff",x"87"),
  1626 => (x"97",x"49",x"a5",x"c2"),
  1627 => (x"a3",x"71",x"4b",x"6c"),
  1628 => (x"4b",x"6b",x"97",x"4b"),
  1629 => (x"6e",x"7e",x"6c",x"97"),
  1630 => (x"c8",x"80",x"c1",x"48"),
  1631 => (x"98",x"c7",x"58",x"a6"),
  1632 => (x"70",x"58",x"a6",x"cc"),
  1633 => (x"e1",x"fe",x"7c",x"97"),
  1634 => (x"f4",x"48",x"73",x"87"),
  1635 => (x"26",x"4d",x"26",x"8e"),
  1636 => (x"26",x"4b",x"26",x"4c"),
  1637 => (x"5b",x"5e",x"0e",x"4f"),
  1638 => (x"86",x"f4",x"0e",x"5c"),
  1639 => (x"66",x"d8",x"4c",x"71"),
  1640 => (x"9a",x"ff",x"c3",x"4a"),
  1641 => (x"97",x"4b",x"a4",x"c2"),
  1642 => (x"a1",x"73",x"49",x"6c"),
  1643 => (x"97",x"51",x"72",x"49"),
  1644 => (x"48",x"6e",x"7e",x"6c"),
  1645 => (x"a6",x"c8",x"80",x"c1"),
  1646 => (x"cc",x"98",x"c7",x"58"),
  1647 => (x"54",x"70",x"58",x"a6"),
  1648 => (x"ca",x"ff",x"8e",x"f4"),
  1649 => (x"fd",x"1e",x"1e",x"87"),
  1650 => (x"bf",x"e0",x"87",x"e8"),
  1651 => (x"e0",x"c0",x"49",x"4a"),
  1652 => (x"cb",x"02",x"99",x"c0"),
  1653 => (x"c2",x"1e",x"72",x"87"),
  1654 => (x"fe",x"49",x"cf",x"f7"),
  1655 => (x"86",x"c4",x"87",x"f7"),
  1656 => (x"70",x"87",x"fd",x"fc"),
  1657 => (x"87",x"c2",x"fd",x"7e"),
  1658 => (x"1e",x"4f",x"26",x"26"),
  1659 => (x"49",x"cf",x"f7",x"c2"),
  1660 => (x"c1",x"87",x"c7",x"fd"),
  1661 => (x"fc",x"49",x"c5",x"e7"),
  1662 => (x"d9",x"c5",x"87",x"da"),
  1663 => (x"0e",x"4f",x"26",x"87"),
  1664 => (x"5d",x"5c",x"5b",x"5e"),
  1665 => (x"ee",x"f7",x"c2",x"0e"),
  1666 => (x"e9",x"c1",x"4a",x"bf"),
  1667 => (x"4c",x"49",x"bf",x"d3"),
  1668 => (x"4d",x"71",x"bc",x"72"),
  1669 => (x"c0",x"87",x"db",x"fc"),
  1670 => (x"d0",x"49",x"74",x"4b"),
  1671 => (x"87",x"d5",x"02",x"99"),
  1672 => (x"99",x"d0",x"49",x"75"),
  1673 => (x"1e",x"c0",x"1e",x"71"),
  1674 => (x"4a",x"e5",x"ef",x"c1"),
  1675 => (x"49",x"12",x"82",x"73"),
  1676 => (x"c8",x"87",x"e4",x"c0"),
  1677 => (x"2d",x"2c",x"c1",x"86"),
  1678 => (x"04",x"ab",x"c8",x"83"),
  1679 => (x"fb",x"87",x"da",x"ff"),
  1680 => (x"e9",x"c1",x"87",x"e8"),
  1681 => (x"f7",x"c2",x"48",x"d3"),
  1682 => (x"26",x"78",x"bf",x"ee"),
  1683 => (x"26",x"4c",x"26",x"4d"),
  1684 => (x"00",x"4f",x"26",x"4b"),
  1685 => (x"1e",x"00",x"00",x"00"),
  1686 => (x"c8",x"48",x"d0",x"ff"),
  1687 => (x"d4",x"ff",x"78",x"e1"),
  1688 => (x"c4",x"78",x"c5",x"48"),
  1689 => (x"87",x"c3",x"02",x"66"),
  1690 => (x"c8",x"78",x"e0",x"c3"),
  1691 => (x"87",x"c6",x"02",x"66"),
  1692 => (x"c3",x"48",x"d4",x"ff"),
  1693 => (x"d4",x"ff",x"78",x"f0"),
  1694 => (x"ff",x"78",x"71",x"48"),
  1695 => (x"e1",x"c8",x"48",x"d0"),
  1696 => (x"78",x"e0",x"c0",x"78"),
  1697 => (x"5e",x"0e",x"4f",x"26"),
  1698 => (x"71",x"0e",x"5c",x"5b"),
  1699 => (x"cf",x"f7",x"c2",x"4c"),
  1700 => (x"87",x"ee",x"fa",x"49"),
  1701 => (x"b7",x"c0",x"4a",x"70"),
  1702 => (x"e3",x"c2",x"04",x"aa"),
  1703 => (x"aa",x"e0",x"c3",x"87"),
  1704 => (x"c1",x"87",x"c9",x"05"),
  1705 => (x"c1",x"48",x"c9",x"ed"),
  1706 => (x"87",x"d4",x"c2",x"78"),
  1707 => (x"05",x"aa",x"f0",x"c3"),
  1708 => (x"ed",x"c1",x"87",x"c9"),
  1709 => (x"78",x"c1",x"48",x"c5"),
  1710 => (x"c1",x"87",x"f5",x"c1"),
  1711 => (x"02",x"bf",x"c9",x"ed"),
  1712 => (x"4b",x"72",x"87",x"c7"),
  1713 => (x"c2",x"b3",x"c0",x"c2"),
  1714 => (x"74",x"4b",x"72",x"87"),
  1715 => (x"87",x"d1",x"05",x"9c"),
  1716 => (x"bf",x"c5",x"ed",x"c1"),
  1717 => (x"c9",x"ed",x"c1",x"1e"),
  1718 => (x"49",x"72",x"1e",x"bf"),
  1719 => (x"c8",x"87",x"f8",x"fd"),
  1720 => (x"c5",x"ed",x"c1",x"86"),
  1721 => (x"e0",x"c0",x"02",x"bf"),
  1722 => (x"c4",x"49",x"73",x"87"),
  1723 => (x"c1",x"91",x"29",x"b7"),
  1724 => (x"73",x"81",x"e5",x"ee"),
  1725 => (x"c2",x"9a",x"cf",x"4a"),
  1726 => (x"72",x"48",x"c1",x"92"),
  1727 => (x"ff",x"4a",x"70",x"30"),
  1728 => (x"69",x"48",x"72",x"ba"),
  1729 => (x"db",x"79",x"70",x"98"),
  1730 => (x"c4",x"49",x"73",x"87"),
  1731 => (x"c1",x"91",x"29",x"b7"),
  1732 => (x"73",x"81",x"e5",x"ee"),
  1733 => (x"c2",x"9a",x"cf",x"4a"),
  1734 => (x"72",x"48",x"c3",x"92"),
  1735 => (x"48",x"4a",x"70",x"30"),
  1736 => (x"79",x"70",x"b0",x"69"),
  1737 => (x"48",x"c9",x"ed",x"c1"),
  1738 => (x"ed",x"c1",x"78",x"c0"),
  1739 => (x"78",x"c0",x"48",x"c5"),
  1740 => (x"49",x"cf",x"f7",x"c2"),
  1741 => (x"70",x"87",x"cb",x"f8"),
  1742 => (x"aa",x"b7",x"c0",x"4a"),
  1743 => (x"87",x"dd",x"fd",x"03"),
  1744 => (x"c8",x"fc",x"48",x"c0"),
  1745 => (x"00",x"00",x"00",x"87"),
  1746 => (x"00",x"00",x"00",x"00"),
  1747 => (x"4a",x"71",x"1e",x"00"),
  1748 => (x"87",x"f2",x"fc",x"49"),
  1749 => (x"c0",x"1e",x"4f",x"26"),
  1750 => (x"c4",x"49",x"72",x"4a"),
  1751 => (x"e5",x"ee",x"c1",x"91"),
  1752 => (x"c1",x"79",x"c0",x"81"),
  1753 => (x"aa",x"b7",x"d0",x"82"),
  1754 => (x"26",x"87",x"ee",x"04"),
  1755 => (x"5b",x"5e",x"0e",x"4f"),
  1756 => (x"71",x"0e",x"5d",x"5c"),
  1757 => (x"87",x"fa",x"f6",x"4d"),
  1758 => (x"b7",x"c4",x"4a",x"75"),
  1759 => (x"ee",x"c1",x"92",x"2a"),
  1760 => (x"4c",x"75",x"82",x"e5"),
  1761 => (x"94",x"c2",x"9c",x"cf"),
  1762 => (x"74",x"4b",x"49",x"6a"),
  1763 => (x"c2",x"9b",x"c3",x"2b"),
  1764 => (x"70",x"30",x"74",x"48"),
  1765 => (x"74",x"bc",x"ff",x"4c"),
  1766 => (x"70",x"98",x"71",x"48"),
  1767 => (x"87",x"ca",x"f6",x"7a"),
  1768 => (x"e6",x"fa",x"48",x"73"),
  1769 => (x"00",x"00",x"00",x"87"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"26",x"1e",x"16",x"00"),
  1786 => (x"3d",x"36",x"2e",x"25"),
  1787 => (x"d0",x"ff",x"1e",x"3e"),
  1788 => (x"78",x"e1",x"c8",x"48"),
  1789 => (x"d4",x"ff",x"48",x"71"),
  1790 => (x"4f",x"26",x"78",x"08"),
  1791 => (x"48",x"d0",x"ff",x"1e"),
  1792 => (x"71",x"78",x"e1",x"c8"),
  1793 => (x"08",x"d4",x"ff",x"48"),
  1794 => (x"48",x"66",x"c4",x"78"),
  1795 => (x"78",x"08",x"d4",x"ff"),
  1796 => (x"71",x"1e",x"4f",x"26"),
  1797 => (x"49",x"66",x"c4",x"4a"),
  1798 => (x"ff",x"49",x"72",x"1e"),
  1799 => (x"d0",x"ff",x"87",x"de"),
  1800 => (x"78",x"e0",x"c0",x"48"),
  1801 => (x"1e",x"4f",x"26",x"26"),
  1802 => (x"b7",x"c2",x"4a",x"71"),
  1803 => (x"87",x"c3",x"03",x"aa"),
  1804 => (x"ce",x"87",x"c2",x"82"),
  1805 => (x"1e",x"66",x"c4",x"82"),
  1806 => (x"d5",x"ff",x"49",x"72"),
  1807 => (x"4f",x"26",x"26",x"87"),
  1808 => (x"4a",x"d4",x"ff",x"1e"),
  1809 => (x"ff",x"7a",x"ff",x"c3"),
  1810 => (x"e1",x"c8",x"48",x"d0"),
  1811 => (x"c2",x"7a",x"de",x"78"),
  1812 => (x"7a",x"bf",x"d9",x"f7"),
  1813 => (x"28",x"c8",x"48",x"49"),
  1814 => (x"48",x"71",x"7a",x"70"),
  1815 => (x"7a",x"70",x"28",x"d0"),
  1816 => (x"28",x"d8",x"48",x"71"),
  1817 => (x"d0",x"ff",x"7a",x"70"),
  1818 => (x"78",x"e0",x"c0",x"48"),
  1819 => (x"5e",x"0e",x"4f",x"26"),
  1820 => (x"0e",x"5d",x"5c",x"5b"),
  1821 => (x"f7",x"c2",x"4c",x"71"),
  1822 => (x"4b",x"4d",x"bf",x"d9"),
  1823 => (x"66",x"d0",x"2b",x"74"),
  1824 => (x"d4",x"83",x"c1",x"9b"),
  1825 => (x"c2",x"04",x"ab",x"66"),
  1826 => (x"74",x"4b",x"c0",x"87"),
  1827 => (x"49",x"66",x"d0",x"4a"),
  1828 => (x"b9",x"ff",x"31",x"72"),
  1829 => (x"48",x"73",x"99",x"75"),
  1830 => (x"4a",x"70",x"30",x"72"),
  1831 => (x"c2",x"b0",x"71",x"48"),
  1832 => (x"fe",x"58",x"dd",x"f7"),
  1833 => (x"4d",x"26",x"87",x"da"),
  1834 => (x"4b",x"26",x"4c",x"26"),
  1835 => (x"ff",x"1e",x"4f",x"26"),
  1836 => (x"c9",x"c8",x"48",x"d0"),
  1837 => (x"ff",x"48",x"71",x"78"),
  1838 => (x"26",x"78",x"08",x"d4"),
  1839 => (x"4a",x"71",x"1e",x"4f"),
  1840 => (x"ff",x"87",x"eb",x"49"),
  1841 => (x"78",x"c8",x"48",x"d0"),
  1842 => (x"73",x"1e",x"4f",x"26"),
  1843 => (x"c2",x"4b",x"71",x"1e"),
  1844 => (x"02",x"bf",x"e9",x"f7"),
  1845 => (x"eb",x"c2",x"87",x"c3"),
  1846 => (x"48",x"d0",x"ff",x"87"),
  1847 => (x"73",x"78",x"c9",x"c8"),
  1848 => (x"b1",x"e0",x"c0",x"49"),
  1849 => (x"71",x"48",x"d4",x"ff"),
  1850 => (x"dd",x"f7",x"c2",x"78"),
  1851 => (x"c8",x"78",x"c0",x"48"),
  1852 => (x"87",x"c5",x"02",x"66"),
  1853 => (x"c2",x"49",x"ff",x"c3"),
  1854 => (x"c2",x"49",x"c0",x"87"),
  1855 => (x"cc",x"59",x"e5",x"f7"),
  1856 => (x"87",x"c6",x"02",x"66"),
  1857 => (x"4a",x"d5",x"d5",x"c5"),
  1858 => (x"ff",x"cf",x"87",x"c4"),
  1859 => (x"f7",x"c2",x"4a",x"ff"),
  1860 => (x"f7",x"c2",x"5a",x"e9"),
  1861 => (x"78",x"c1",x"48",x"e9"),
  1862 => (x"4d",x"26",x"87",x"c4"),
  1863 => (x"4b",x"26",x"4c",x"26"),
  1864 => (x"5e",x"0e",x"4f",x"26"),
  1865 => (x"0e",x"5d",x"5c",x"5b"),
  1866 => (x"f7",x"c2",x"4a",x"71"),
  1867 => (x"72",x"4c",x"bf",x"e5"),
  1868 => (x"87",x"cb",x"02",x"9a"),
  1869 => (x"c1",x"91",x"c8",x"49"),
  1870 => (x"71",x"4b",x"c0",x"f3"),
  1871 => (x"c1",x"87",x"c4",x"83"),
  1872 => (x"c0",x"4b",x"c0",x"f7"),
  1873 => (x"74",x"49",x"13",x"4d"),
  1874 => (x"e1",x"f7",x"c2",x"99"),
  1875 => (x"d4",x"ff",x"b9",x"bf"),
  1876 => (x"c1",x"78",x"71",x"48"),
  1877 => (x"c8",x"85",x"2c",x"b7"),
  1878 => (x"e8",x"04",x"ad",x"b7"),
  1879 => (x"dd",x"f7",x"c2",x"87"),
  1880 => (x"80",x"c8",x"48",x"bf"),
  1881 => (x"58",x"e1",x"f7",x"c2"),
  1882 => (x"1e",x"87",x"ef",x"fe"),
  1883 => (x"4b",x"71",x"1e",x"73"),
  1884 => (x"02",x"9a",x"4a",x"13"),
  1885 => (x"49",x"72",x"87",x"cb"),
  1886 => (x"13",x"87",x"e7",x"fe"),
  1887 => (x"f5",x"05",x"9a",x"4a"),
  1888 => (x"87",x"da",x"fe",x"87"),
  1889 => (x"dd",x"f7",x"c2",x"1e"),
  1890 => (x"f7",x"c2",x"49",x"bf"),
  1891 => (x"a1",x"c1",x"48",x"dd"),
  1892 => (x"b7",x"c0",x"c4",x"78"),
  1893 => (x"87",x"db",x"03",x"a9"),
  1894 => (x"c2",x"48",x"d4",x"ff"),
  1895 => (x"78",x"bf",x"e1",x"f7"),
  1896 => (x"bf",x"dd",x"f7",x"c2"),
  1897 => (x"dd",x"f7",x"c2",x"49"),
  1898 => (x"78",x"a1",x"c1",x"48"),
  1899 => (x"a9",x"b7",x"c0",x"c4"),
  1900 => (x"ff",x"87",x"e5",x"04"),
  1901 => (x"78",x"c8",x"48",x"d0"),
  1902 => (x"48",x"e9",x"f7",x"c2"),
  1903 => (x"4f",x"26",x"78",x"c0"),
  1904 => (x"00",x"00",x"00",x"00"),
  1905 => (x"00",x"00",x"00",x"00"),
  1906 => (x"5f",x"00",x"00",x"00"),
  1907 => (x"00",x"00",x"00",x"5f"),
  1908 => (x"00",x"03",x"03",x"00"),
  1909 => (x"00",x"00",x"03",x"03"),
  1910 => (x"14",x"7f",x"7f",x"14"),
  1911 => (x"00",x"14",x"7f",x"7f"),
  1912 => (x"6b",x"2e",x"24",x"00"),
  1913 => (x"00",x"12",x"3a",x"6b"),
  1914 => (x"18",x"36",x"6a",x"4c"),
  1915 => (x"00",x"32",x"56",x"6c"),
  1916 => (x"59",x"4f",x"7e",x"30"),
  1917 => (x"40",x"68",x"3a",x"77"),
  1918 => (x"07",x"04",x"00",x"00"),
  1919 => (x"00",x"00",x"00",x"03"),
  1920 => (x"3e",x"1c",x"00",x"00"),
  1921 => (x"00",x"00",x"41",x"63"),
  1922 => (x"63",x"41",x"00",x"00"),
  1923 => (x"00",x"00",x"1c",x"3e"),
  1924 => (x"1c",x"3e",x"2a",x"08"),
  1925 => (x"08",x"2a",x"3e",x"1c"),
  1926 => (x"3e",x"08",x"08",x"00"),
  1927 => (x"00",x"08",x"08",x"3e"),
  1928 => (x"e0",x"80",x"00",x"00"),
  1929 => (x"00",x"00",x"00",x"60"),
  1930 => (x"08",x"08",x"08",x"00"),
  1931 => (x"00",x"08",x"08",x"08"),
  1932 => (x"60",x"00",x"00",x"00"),
  1933 => (x"00",x"00",x"00",x"60"),
  1934 => (x"18",x"30",x"60",x"40"),
  1935 => (x"01",x"03",x"06",x"0c"),
  1936 => (x"59",x"7f",x"3e",x"00"),
  1937 => (x"00",x"3e",x"7f",x"4d"),
  1938 => (x"7f",x"06",x"04",x"00"),
  1939 => (x"00",x"00",x"00",x"7f"),
  1940 => (x"71",x"63",x"42",x"00"),
  1941 => (x"00",x"46",x"4f",x"59"),
  1942 => (x"49",x"63",x"22",x"00"),
  1943 => (x"00",x"36",x"7f",x"49"),
  1944 => (x"13",x"16",x"1c",x"18"),
  1945 => (x"00",x"10",x"7f",x"7f"),
  1946 => (x"45",x"67",x"27",x"00"),
  1947 => (x"00",x"39",x"7d",x"45"),
  1948 => (x"4b",x"7e",x"3c",x"00"),
  1949 => (x"00",x"30",x"79",x"49"),
  1950 => (x"71",x"01",x"01",x"00"),
  1951 => (x"00",x"07",x"0f",x"79"),
  1952 => (x"49",x"7f",x"36",x"00"),
  1953 => (x"00",x"36",x"7f",x"49"),
  1954 => (x"49",x"4f",x"06",x"00"),
  1955 => (x"00",x"1e",x"3f",x"69"),
  1956 => (x"66",x"00",x"00",x"00"),
  1957 => (x"00",x"00",x"00",x"66"),
  1958 => (x"e6",x"80",x"00",x"00"),
  1959 => (x"00",x"00",x"00",x"66"),
  1960 => (x"14",x"08",x"08",x"00"),
  1961 => (x"00",x"22",x"22",x"14"),
  1962 => (x"14",x"14",x"14",x"00"),
  1963 => (x"00",x"14",x"14",x"14"),
  1964 => (x"14",x"22",x"22",x"00"),
  1965 => (x"00",x"08",x"08",x"14"),
  1966 => (x"51",x"03",x"02",x"00"),
  1967 => (x"00",x"06",x"0f",x"59"),
  1968 => (x"5d",x"41",x"7f",x"3e"),
  1969 => (x"00",x"1e",x"1f",x"55"),
  1970 => (x"09",x"7f",x"7e",x"00"),
  1971 => (x"00",x"7e",x"7f",x"09"),
  1972 => (x"49",x"7f",x"7f",x"00"),
  1973 => (x"00",x"36",x"7f",x"49"),
  1974 => (x"63",x"3e",x"1c",x"00"),
  1975 => (x"00",x"41",x"41",x"41"),
  1976 => (x"41",x"7f",x"7f",x"00"),
  1977 => (x"00",x"1c",x"3e",x"63"),
  1978 => (x"49",x"7f",x"7f",x"00"),
  1979 => (x"00",x"41",x"41",x"49"),
  1980 => (x"09",x"7f",x"7f",x"00"),
  1981 => (x"00",x"01",x"01",x"09"),
  1982 => (x"41",x"7f",x"3e",x"00"),
  1983 => (x"00",x"7a",x"7b",x"49"),
  1984 => (x"08",x"7f",x"7f",x"00"),
  1985 => (x"00",x"7f",x"7f",x"08"),
  1986 => (x"7f",x"41",x"00",x"00"),
  1987 => (x"00",x"00",x"41",x"7f"),
  1988 => (x"40",x"60",x"20",x"00"),
  1989 => (x"00",x"3f",x"7f",x"40"),
  1990 => (x"1c",x"08",x"7f",x"7f"),
  1991 => (x"00",x"41",x"63",x"36"),
  1992 => (x"40",x"7f",x"7f",x"00"),
  1993 => (x"00",x"40",x"40",x"40"),
  1994 => (x"0c",x"06",x"7f",x"7f"),
  1995 => (x"00",x"7f",x"7f",x"06"),
  1996 => (x"0c",x"06",x"7f",x"7f"),
  1997 => (x"00",x"7f",x"7f",x"18"),
  1998 => (x"41",x"7f",x"3e",x"00"),
  1999 => (x"00",x"3e",x"7f",x"41"),
  2000 => (x"09",x"7f",x"7f",x"00"),
  2001 => (x"00",x"06",x"0f",x"09"),
  2002 => (x"61",x"41",x"7f",x"3e"),
  2003 => (x"00",x"40",x"7e",x"7f"),
  2004 => (x"09",x"7f",x"7f",x"00"),
  2005 => (x"00",x"66",x"7f",x"19"),
  2006 => (x"4d",x"6f",x"26",x"00"),
  2007 => (x"00",x"32",x"7b",x"59"),
  2008 => (x"7f",x"01",x"01",x"00"),
  2009 => (x"00",x"01",x"01",x"7f"),
  2010 => (x"40",x"7f",x"3f",x"00"),
  2011 => (x"00",x"3f",x"7f",x"40"),
  2012 => (x"70",x"3f",x"0f",x"00"),
  2013 => (x"00",x"0f",x"3f",x"70"),
  2014 => (x"18",x"30",x"7f",x"7f"),
  2015 => (x"00",x"7f",x"7f",x"30"),
  2016 => (x"1c",x"36",x"63",x"41"),
  2017 => (x"41",x"63",x"36",x"1c"),
  2018 => (x"7c",x"06",x"03",x"01"),
  2019 => (x"01",x"03",x"06",x"7c"),
  2020 => (x"4d",x"59",x"71",x"61"),
  2021 => (x"00",x"41",x"43",x"47"),
  2022 => (x"7f",x"7f",x"00",x"00"),
  2023 => (x"00",x"00",x"41",x"41"),
  2024 => (x"0c",x"06",x"03",x"01"),
  2025 => (x"40",x"60",x"30",x"18"),
  2026 => (x"41",x"41",x"00",x"00"),
  2027 => (x"00",x"00",x"7f",x"7f"),
  2028 => (x"03",x"06",x"0c",x"08"),
  2029 => (x"00",x"08",x"0c",x"06"),
  2030 => (x"80",x"80",x"80",x"80"),
  2031 => (x"00",x"80",x"80",x"80"),
  2032 => (x"03",x"00",x"00",x"00"),
  2033 => (x"00",x"00",x"04",x"07"),
  2034 => (x"54",x"74",x"20",x"00"),
  2035 => (x"00",x"78",x"7c",x"54"),
  2036 => (x"44",x"7f",x"7f",x"00"),
  2037 => (x"00",x"38",x"7c",x"44"),
  2038 => (x"44",x"7c",x"38",x"00"),
  2039 => (x"00",x"00",x"44",x"44"),
  2040 => (x"44",x"7c",x"38",x"00"),
  2041 => (x"00",x"7f",x"7f",x"44"),
  2042 => (x"54",x"7c",x"38",x"00"),
  2043 => (x"00",x"18",x"5c",x"54"),
  2044 => (x"7f",x"7e",x"04",x"00"),
  2045 => (x"00",x"00",x"05",x"05"),
  2046 => (x"a4",x"bc",x"18",x"00"),
  2047 => (x"00",x"7c",x"fc",x"a4"),
  2048 => (x"04",x"7f",x"7f",x"00"),
  2049 => (x"00",x"78",x"7c",x"04"),
  2050 => (x"3d",x"00",x"00",x"00"),
  2051 => (x"00",x"00",x"40",x"7d"),
  2052 => (x"80",x"80",x"80",x"00"),
  2053 => (x"00",x"00",x"7d",x"fd"),
  2054 => (x"10",x"7f",x"7f",x"00"),
  2055 => (x"00",x"44",x"6c",x"38"),
  2056 => (x"3f",x"00",x"00",x"00"),
  2057 => (x"00",x"00",x"40",x"7f"),
  2058 => (x"18",x"0c",x"7c",x"7c"),
  2059 => (x"00",x"78",x"7c",x"0c"),
  2060 => (x"04",x"7c",x"7c",x"00"),
  2061 => (x"00",x"78",x"7c",x"04"),
  2062 => (x"44",x"7c",x"38",x"00"),
  2063 => (x"00",x"38",x"7c",x"44"),
  2064 => (x"24",x"fc",x"fc",x"00"),
  2065 => (x"00",x"18",x"3c",x"24"),
  2066 => (x"24",x"3c",x"18",x"00"),
  2067 => (x"00",x"fc",x"fc",x"24"),
  2068 => (x"04",x"7c",x"7c",x"00"),
  2069 => (x"00",x"08",x"0c",x"04"),
  2070 => (x"54",x"5c",x"48",x"00"),
  2071 => (x"00",x"20",x"74",x"54"),
  2072 => (x"7f",x"3f",x"04",x"00"),
  2073 => (x"00",x"00",x"44",x"44"),
  2074 => (x"40",x"7c",x"3c",x"00"),
  2075 => (x"00",x"7c",x"7c",x"40"),
  2076 => (x"60",x"3c",x"1c",x"00"),
  2077 => (x"00",x"1c",x"3c",x"60"),
  2078 => (x"30",x"60",x"7c",x"3c"),
  2079 => (x"00",x"3c",x"7c",x"60"),
  2080 => (x"10",x"38",x"6c",x"44"),
  2081 => (x"00",x"44",x"6c",x"38"),
  2082 => (x"e0",x"bc",x"1c",x"00"),
  2083 => (x"00",x"1c",x"3c",x"60"),
  2084 => (x"74",x"64",x"44",x"00"),
  2085 => (x"00",x"44",x"4c",x"5c"),
  2086 => (x"3e",x"08",x"08",x"00"),
  2087 => (x"00",x"41",x"41",x"77"),
  2088 => (x"7f",x"00",x"00",x"00"),
  2089 => (x"00",x"00",x"00",x"7f"),
  2090 => (x"77",x"41",x"41",x"00"),
  2091 => (x"00",x"08",x"08",x"3e"),
  2092 => (x"03",x"01",x"01",x"02"),
  2093 => (x"00",x"01",x"02",x"02"),
  2094 => (x"7f",x"7f",x"7f",x"7f"),
  2095 => (x"00",x"7f",x"7f",x"7f"),
  2096 => (x"1c",x"1c",x"08",x"08"),
  2097 => (x"7f",x"7f",x"3e",x"3e"),
  2098 => (x"3e",x"3e",x"7f",x"7f"),
  2099 => (x"08",x"08",x"1c",x"1c"),
  2100 => (x"7c",x"18",x"10",x"00"),
  2101 => (x"00",x"10",x"18",x"7c"),
  2102 => (x"7c",x"30",x"10",x"00"),
  2103 => (x"00",x"10",x"30",x"7c"),
  2104 => (x"60",x"60",x"30",x"10"),
  2105 => (x"00",x"06",x"1e",x"78"),
  2106 => (x"18",x"3c",x"66",x"42"),
  2107 => (x"00",x"42",x"66",x"3c"),
  2108 => (x"c2",x"6a",x"38",x"78"),
  2109 => (x"00",x"38",x"6c",x"c6"),
  2110 => (x"60",x"00",x"00",x"60"),
  2111 => (x"00",x"60",x"00",x"00"),
  2112 => (x"5c",x"5b",x"5e",x"0e"),
  2113 => (x"71",x"1e",x"0e",x"5d"),
  2114 => (x"fa",x"f7",x"c2",x"4c"),
  2115 => (x"4b",x"c0",x"4d",x"bf"),
  2116 => (x"ab",x"74",x"1e",x"c0"),
  2117 => (x"c4",x"87",x"c7",x"02"),
  2118 => (x"78",x"c0",x"48",x"a6"),
  2119 => (x"a6",x"c4",x"87",x"c5"),
  2120 => (x"c4",x"78",x"c1",x"48"),
  2121 => (x"49",x"73",x"1e",x"66"),
  2122 => (x"c8",x"87",x"df",x"ee"),
  2123 => (x"49",x"e0",x"c0",x"86"),
  2124 => (x"c4",x"87",x"ef",x"ef"),
  2125 => (x"49",x"6a",x"4a",x"a5"),
  2126 => (x"f1",x"87",x"f0",x"f0"),
  2127 => (x"85",x"cb",x"87",x"c6"),
  2128 => (x"b7",x"c8",x"83",x"c1"),
  2129 => (x"c7",x"ff",x"04",x"ab"),
  2130 => (x"4d",x"26",x"26",x"87"),
  2131 => (x"4b",x"26",x"4c",x"26"),
  2132 => (x"71",x"1e",x"4f",x"26"),
  2133 => (x"fe",x"f7",x"c2",x"4a"),
  2134 => (x"fe",x"f7",x"c2",x"5a"),
  2135 => (x"49",x"78",x"c7",x"48"),
  2136 => (x"26",x"87",x"dd",x"fe"),
  2137 => (x"1e",x"73",x"1e",x"4f"),
  2138 => (x"b7",x"c0",x"4a",x"71"),
  2139 => (x"87",x"d3",x"03",x"aa"),
  2140 => (x"bf",x"f2",x"d5",x"c2"),
  2141 => (x"c1",x"87",x"c4",x"05"),
  2142 => (x"c0",x"87",x"c2",x"4b"),
  2143 => (x"f6",x"d5",x"c2",x"4b"),
  2144 => (x"c2",x"87",x"c4",x"5b"),
  2145 => (x"c2",x"5a",x"f6",x"d5"),
  2146 => (x"4a",x"bf",x"f2",x"d5"),
  2147 => (x"c0",x"c1",x"9a",x"c1"),
  2148 => (x"e8",x"ec",x"49",x"a2"),
  2149 => (x"da",x"d5",x"c2",x"87"),
  2150 => (x"d5",x"c2",x"49",x"bf"),
  2151 => (x"fc",x"b1",x"bf",x"f2"),
  2152 => (x"fe",x"78",x"71",x"48"),
  2153 => (x"71",x"1e",x"87",x"e8"),
  2154 => (x"1e",x"66",x"c4",x"4a"),
  2155 => (x"f6",x"e9",x"49",x"72"),
  2156 => (x"4f",x"26",x"26",x"87"),
  2157 => (x"f2",x"d5",x"c2",x"1e"),
  2158 => (x"d0",x"e6",x"49",x"bf"),
  2159 => (x"f2",x"f7",x"c2",x"87"),
  2160 => (x"78",x"bf",x"e8",x"48"),
  2161 => (x"48",x"ee",x"f7",x"c2"),
  2162 => (x"c2",x"78",x"bf",x"ec"),
  2163 => (x"4a",x"bf",x"f2",x"f7"),
  2164 => (x"99",x"ff",x"c3",x"49"),
  2165 => (x"72",x"2a",x"b7",x"c8"),
  2166 => (x"c2",x"b0",x"71",x"48"),
  2167 => (x"26",x"58",x"fa",x"f7"),
  2168 => (x"5b",x"5e",x"0e",x"4f"),
  2169 => (x"71",x"0e",x"5d",x"5c"),
  2170 => (x"87",x"c8",x"ff",x"4b"),
  2171 => (x"48",x"ed",x"f7",x"c2"),
  2172 => (x"49",x"73",x"50",x"c0"),
  2173 => (x"70",x"87",x"f6",x"e5"),
  2174 => (x"9c",x"c2",x"4c",x"49"),
  2175 => (x"cd",x"49",x"ee",x"cb"),
  2176 => (x"49",x"70",x"87",x"f8"),
  2177 => (x"ed",x"f7",x"c2",x"4d"),
  2178 => (x"c1",x"05",x"bf",x"97"),
  2179 => (x"66",x"d0",x"87",x"e2"),
  2180 => (x"f6",x"f7",x"c2",x"49"),
  2181 => (x"d6",x"05",x"99",x"bf"),
  2182 => (x"49",x"66",x"d4",x"87"),
  2183 => (x"bf",x"ee",x"f7",x"c2"),
  2184 => (x"87",x"cb",x"05",x"99"),
  2185 => (x"c4",x"e5",x"49",x"73"),
  2186 => (x"02",x"98",x"70",x"87"),
  2187 => (x"c1",x"87",x"c1",x"c1"),
  2188 => (x"87",x"c0",x"fe",x"4c"),
  2189 => (x"cd",x"cd",x"49",x"75"),
  2190 => (x"02",x"98",x"70",x"87"),
  2191 => (x"f7",x"c2",x"87",x"c6"),
  2192 => (x"50",x"c1",x"48",x"ed"),
  2193 => (x"97",x"ed",x"f7",x"c2"),
  2194 => (x"e3",x"c0",x"05",x"bf"),
  2195 => (x"f6",x"f7",x"c2",x"87"),
  2196 => (x"66",x"d0",x"49",x"bf"),
  2197 => (x"d6",x"ff",x"05",x"99"),
  2198 => (x"ee",x"f7",x"c2",x"87"),
  2199 => (x"66",x"d4",x"49",x"bf"),
  2200 => (x"ca",x"ff",x"05",x"99"),
  2201 => (x"e4",x"49",x"73",x"87"),
  2202 => (x"98",x"70",x"87",x"c3"),
  2203 => (x"87",x"ff",x"fe",x"05"),
  2204 => (x"d5",x"fb",x"48",x"74"),
  2205 => (x"5b",x"5e",x"0e",x"87"),
  2206 => (x"f8",x"0e",x"5d",x"5c"),
  2207 => (x"4c",x"4d",x"c0",x"86"),
  2208 => (x"c4",x"7e",x"bf",x"ec"),
  2209 => (x"f7",x"c2",x"48",x"a6"),
  2210 => (x"c0",x"78",x"bf",x"fa"),
  2211 => (x"f7",x"c1",x"1e",x"1e"),
  2212 => (x"87",x"cd",x"fd",x"49"),
  2213 => (x"98",x"70",x"86",x"c8"),
  2214 => (x"87",x"f3",x"c0",x"02"),
  2215 => (x"bf",x"da",x"d5",x"c2"),
  2216 => (x"c1",x"87",x"c4",x"05"),
  2217 => (x"c0",x"87",x"c2",x"7e"),
  2218 => (x"da",x"d5",x"c2",x"7e"),
  2219 => (x"ca",x"78",x"6e",x"48"),
  2220 => (x"66",x"c4",x"1e",x"fc"),
  2221 => (x"c4",x"87",x"c9",x"02"),
  2222 => (x"d3",x"c2",x"48",x"a6"),
  2223 => (x"87",x"c7",x"78",x"f1"),
  2224 => (x"c2",x"48",x"a6",x"c4"),
  2225 => (x"c4",x"78",x"fc",x"d3"),
  2226 => (x"fb",x"c8",x"49",x"66"),
  2227 => (x"c1",x"86",x"c4",x"87"),
  2228 => (x"c7",x"1e",x"c0",x"1e"),
  2229 => (x"87",x"c9",x"fc",x"49"),
  2230 => (x"98",x"70",x"86",x"c8"),
  2231 => (x"ff",x"87",x"cd",x"02"),
  2232 => (x"87",x"c1",x"fa",x"49"),
  2233 => (x"e2",x"49",x"da",x"c1"),
  2234 => (x"4d",x"c1",x"87",x"c3"),
  2235 => (x"97",x"ed",x"f7",x"c2"),
  2236 => (x"87",x"c3",x"02",x"bf"),
  2237 => (x"c2",x"87",x"cd",x"d7"),
  2238 => (x"4b",x"bf",x"f2",x"f7"),
  2239 => (x"bf",x"f2",x"d5",x"c2"),
  2240 => (x"87",x"e1",x"c1",x"05"),
  2241 => (x"bf",x"da",x"d5",x"c2"),
  2242 => (x"87",x"f0",x"c0",x"02"),
  2243 => (x"c8",x"48",x"a6",x"c4"),
  2244 => (x"c2",x"78",x"c0",x"c0"),
  2245 => (x"6e",x"7e",x"de",x"d5"),
  2246 => (x"6e",x"49",x"bf",x"97"),
  2247 => (x"70",x"80",x"c1",x"48"),
  2248 => (x"c8",x"e1",x"71",x"7e"),
  2249 => (x"02",x"98",x"70",x"87"),
  2250 => (x"66",x"c4",x"87",x"c3"),
  2251 => (x"48",x"66",x"c4",x"b3"),
  2252 => (x"c8",x"28",x"b7",x"c1"),
  2253 => (x"98",x"70",x"58",x"a6"),
  2254 => (x"87",x"db",x"ff",x"05"),
  2255 => (x"e0",x"49",x"fd",x"c3"),
  2256 => (x"fa",x"c3",x"87",x"eb"),
  2257 => (x"87",x"e5",x"e0",x"49"),
  2258 => (x"ff",x"c3",x"49",x"73"),
  2259 => (x"c0",x"1e",x"71",x"99"),
  2260 => (x"87",x"d2",x"f9",x"49"),
  2261 => (x"b7",x"c8",x"49",x"73"),
  2262 => (x"c1",x"1e",x"71",x"29"),
  2263 => (x"87",x"c6",x"f9",x"49"),
  2264 => (x"c7",x"c6",x"86",x"c8"),
  2265 => (x"f6",x"f7",x"c2",x"87"),
  2266 => (x"02",x"9b",x"4b",x"bf"),
  2267 => (x"d5",x"c2",x"87",x"df"),
  2268 => (x"c8",x"49",x"bf",x"ee"),
  2269 => (x"98",x"70",x"87",x"d0"),
  2270 => (x"87",x"c4",x"c0",x"05"),
  2271 => (x"87",x"d3",x"4b",x"c0"),
  2272 => (x"c7",x"49",x"e0",x"c2"),
  2273 => (x"d5",x"c2",x"87",x"f4"),
  2274 => (x"c6",x"c0",x"58",x"f2"),
  2275 => (x"ee",x"d5",x"c2",x"87"),
  2276 => (x"73",x"78",x"c0",x"48"),
  2277 => (x"05",x"99",x"c2",x"49"),
  2278 => (x"c3",x"87",x"cf",x"c0"),
  2279 => (x"df",x"ff",x"49",x"eb"),
  2280 => (x"49",x"70",x"87",x"cb"),
  2281 => (x"c0",x"02",x"99",x"c2"),
  2282 => (x"4c",x"fb",x"87",x"c2"),
  2283 => (x"99",x"c1",x"49",x"73"),
  2284 => (x"87",x"cf",x"c0",x"05"),
  2285 => (x"ff",x"49",x"f4",x"c3"),
  2286 => (x"70",x"87",x"f2",x"de"),
  2287 => (x"02",x"99",x"c2",x"49"),
  2288 => (x"fa",x"87",x"c2",x"c0"),
  2289 => (x"c8",x"49",x"73",x"4c"),
  2290 => (x"cf",x"c0",x"05",x"99"),
  2291 => (x"49",x"f5",x"c3",x"87"),
  2292 => (x"87",x"d9",x"de",x"ff"),
  2293 => (x"99",x"c2",x"49",x"70"),
  2294 => (x"87",x"d6",x"c0",x"02"),
  2295 => (x"bf",x"fe",x"f7",x"c2"),
  2296 => (x"87",x"ca",x"c0",x"02"),
  2297 => (x"c2",x"88",x"c1",x"48"),
  2298 => (x"c0",x"58",x"c2",x"f8"),
  2299 => (x"4c",x"ff",x"87",x"c2"),
  2300 => (x"49",x"73",x"4d",x"c1"),
  2301 => (x"c0",x"05",x"99",x"c4"),
  2302 => (x"f2",x"c3",x"87",x"cf"),
  2303 => (x"ec",x"dd",x"ff",x"49"),
  2304 => (x"c2",x"49",x"70",x"87"),
  2305 => (x"dc",x"c0",x"02",x"99"),
  2306 => (x"fe",x"f7",x"c2",x"87"),
  2307 => (x"c7",x"48",x"7e",x"bf"),
  2308 => (x"c0",x"03",x"a8",x"b7"),
  2309 => (x"48",x"6e",x"87",x"cb"),
  2310 => (x"f8",x"c2",x"80",x"c1"),
  2311 => (x"c2",x"c0",x"58",x"c2"),
  2312 => (x"c1",x"4c",x"fe",x"87"),
  2313 => (x"49",x"fd",x"c3",x"4d"),
  2314 => (x"87",x"c1",x"dd",x"ff"),
  2315 => (x"99",x"c2",x"49",x"70"),
  2316 => (x"87",x"d5",x"c0",x"02"),
  2317 => (x"bf",x"fe",x"f7",x"c2"),
  2318 => (x"87",x"c9",x"c0",x"02"),
  2319 => (x"48",x"fe",x"f7",x"c2"),
  2320 => (x"c2",x"c0",x"78",x"c0"),
  2321 => (x"c1",x"4c",x"fd",x"87"),
  2322 => (x"49",x"fa",x"c3",x"4d"),
  2323 => (x"87",x"dd",x"dc",x"ff"),
  2324 => (x"99",x"c2",x"49",x"70"),
  2325 => (x"87",x"d9",x"c0",x"02"),
  2326 => (x"bf",x"fe",x"f7",x"c2"),
  2327 => (x"a8",x"b7",x"c7",x"48"),
  2328 => (x"87",x"c9",x"c0",x"03"),
  2329 => (x"48",x"fe",x"f7",x"c2"),
  2330 => (x"c2",x"c0",x"78",x"c7"),
  2331 => (x"c1",x"4c",x"fc",x"87"),
  2332 => (x"ac",x"b7",x"c0",x"4d"),
  2333 => (x"87",x"d5",x"c0",x"03"),
  2334 => (x"c1",x"48",x"66",x"c4"),
  2335 => (x"7e",x"70",x"80",x"d8"),
  2336 => (x"c0",x"02",x"bf",x"6e"),
  2337 => (x"bf",x"6e",x"87",x"c7"),
  2338 => (x"73",x"49",x"74",x"4b"),
  2339 => (x"c3",x"1e",x"c0",x"0f"),
  2340 => (x"da",x"c1",x"1e",x"f0"),
  2341 => (x"87",x"c9",x"f5",x"49"),
  2342 => (x"98",x"70",x"86",x"c8"),
  2343 => (x"87",x"d9",x"c0",x"02"),
  2344 => (x"bf",x"fe",x"f7",x"c2"),
  2345 => (x"cb",x"49",x"6e",x"7e"),
  2346 => (x"4a",x"66",x"c4",x"91"),
  2347 => (x"02",x"6a",x"82",x"71"),
  2348 => (x"6a",x"87",x"c6",x"c0"),
  2349 => (x"73",x"49",x"6e",x"4b"),
  2350 => (x"02",x"9d",x"75",x"0f"),
  2351 => (x"c2",x"87",x"c8",x"c0"),
  2352 => (x"49",x"bf",x"fe",x"f7"),
  2353 => (x"c2",x"87",x"f9",x"f0"),
  2354 => (x"02",x"bf",x"f6",x"d5"),
  2355 => (x"49",x"87",x"dd",x"c0"),
  2356 => (x"70",x"87",x"f3",x"c2"),
  2357 => (x"d3",x"c0",x"02",x"98"),
  2358 => (x"fe",x"f7",x"c2",x"87"),
  2359 => (x"df",x"f0",x"49",x"bf"),
  2360 => (x"f1",x"49",x"c0",x"87"),
  2361 => (x"d5",x"c2",x"87",x"ff"),
  2362 => (x"78",x"c0",x"48",x"f6"),
  2363 => (x"d9",x"f1",x"8e",x"f8"),
  2364 => (x"79",x"6f",x"4a",x"87"),
  2365 => (x"73",x"79",x"65",x"6b"),
  2366 => (x"00",x"6e",x"6f",x"20"),
  2367 => (x"6b",x"79",x"6f",x"4a"),
  2368 => (x"20",x"73",x"79",x"65"),
  2369 => (x"00",x"66",x"66",x"6f"),
  2370 => (x"5c",x"5b",x"5e",x"0e"),
  2371 => (x"71",x"1e",x"0e",x"5d"),
  2372 => (x"fa",x"f7",x"c2",x"4c"),
  2373 => (x"cd",x"c1",x"49",x"bf"),
  2374 => (x"d1",x"c1",x"4d",x"a1"),
  2375 => (x"74",x"7e",x"69",x"81"),
  2376 => (x"87",x"cf",x"02",x"9c"),
  2377 => (x"74",x"4b",x"a5",x"c4"),
  2378 => (x"fa",x"f7",x"c2",x"7b"),
  2379 => (x"e1",x"f0",x"49",x"bf"),
  2380 => (x"74",x"7b",x"6e",x"87"),
  2381 => (x"87",x"c4",x"05",x"9c"),
  2382 => (x"87",x"c2",x"4b",x"c0"),
  2383 => (x"49",x"73",x"4b",x"c1"),
  2384 => (x"d4",x"87",x"e2",x"f0"),
  2385 => (x"87",x"c8",x"02",x"66"),
  2386 => (x"87",x"ee",x"c0",x"49"),
  2387 => (x"87",x"c2",x"4a",x"70"),
  2388 => (x"d5",x"c2",x"4a",x"c0"),
  2389 => (x"ef",x"26",x"5a",x"fa"),
  2390 => (x"00",x"00",x"87",x"f0"),
  2391 => (x"12",x"58",x"00",x"00"),
  2392 => (x"1b",x"1d",x"14",x"11"),
  2393 => (x"59",x"5a",x"23",x"1c"),
  2394 => (x"f2",x"f5",x"94",x"91"),
  2395 => (x"00",x"00",x"f4",x"eb"),
  2396 => (x"00",x"00",x"00",x"00"),
  2397 => (x"00",x"00",x"00",x"00"),
  2398 => (x"71",x"1e",x"00",x"00"),
  2399 => (x"bf",x"c8",x"ff",x"4a"),
  2400 => (x"48",x"a1",x"72",x"49"),
  2401 => (x"ff",x"1e",x"4f",x"26"),
  2402 => (x"fe",x"89",x"bf",x"c8"),
  2403 => (x"c0",x"c0",x"c0",x"c0"),
  2404 => (x"c4",x"01",x"a9",x"c0"),
  2405 => (x"c2",x"4a",x"c0",x"87"),
  2406 => (x"72",x"4a",x"c1",x"87"),
  2407 => (x"0e",x"4f",x"26",x"48"),
  2408 => (x"5d",x"5c",x"5b",x"5e"),
  2409 => (x"ff",x"4b",x"71",x"0e"),
  2410 => (x"66",x"d0",x"4c",x"d4"),
  2411 => (x"d6",x"78",x"c0",x"48"),
  2412 => (x"f8",x"d8",x"ff",x"49"),
  2413 => (x"7c",x"ff",x"c3",x"87"),
  2414 => (x"ff",x"c3",x"49",x"6c"),
  2415 => (x"49",x"4d",x"71",x"99"),
  2416 => (x"c1",x"99",x"f0",x"c3"),
  2417 => (x"cb",x"05",x"a9",x"e0"),
  2418 => (x"7c",x"ff",x"c3",x"87"),
  2419 => (x"98",x"c3",x"48",x"6c"),
  2420 => (x"78",x"08",x"66",x"d0"),
  2421 => (x"6c",x"7c",x"ff",x"c3"),
  2422 => (x"31",x"c8",x"49",x"4a"),
  2423 => (x"6c",x"7c",x"ff",x"c3"),
  2424 => (x"72",x"b2",x"71",x"4a"),
  2425 => (x"c3",x"31",x"c8",x"49"),
  2426 => (x"4a",x"6c",x"7c",x"ff"),
  2427 => (x"49",x"72",x"b2",x"71"),
  2428 => (x"ff",x"c3",x"31",x"c8"),
  2429 => (x"71",x"4a",x"6c",x"7c"),
  2430 => (x"48",x"d0",x"ff",x"b2"),
  2431 => (x"73",x"78",x"e0",x"c0"),
  2432 => (x"87",x"c2",x"02",x"9b"),
  2433 => (x"48",x"75",x"7b",x"72"),
  2434 => (x"4c",x"26",x"4d",x"26"),
  2435 => (x"4f",x"26",x"4b",x"26"),
  2436 => (x"0e",x"4f",x"26",x"1e"),
  2437 => (x"0e",x"5c",x"5b",x"5e"),
  2438 => (x"1e",x"76",x"86",x"f8"),
  2439 => (x"fd",x"49",x"a6",x"c8"),
  2440 => (x"86",x"c4",x"87",x"fd"),
  2441 => (x"48",x"6e",x"4b",x"70"),
  2442 => (x"c3",x"03",x"a8",x"c2"),
  2443 => (x"4a",x"73",x"87",x"c6"),
  2444 => (x"c1",x"9a",x"f0",x"c3"),
  2445 => (x"c7",x"02",x"aa",x"d0"),
  2446 => (x"aa",x"e0",x"c1",x"87"),
  2447 => (x"87",x"f4",x"c2",x"05"),
  2448 => (x"99",x"c8",x"49",x"73"),
  2449 => (x"ff",x"87",x"c3",x"02"),
  2450 => (x"4c",x"73",x"87",x"c6"),
  2451 => (x"ac",x"c2",x"9c",x"c3"),
  2452 => (x"87",x"cd",x"c1",x"05"),
  2453 => (x"c9",x"49",x"66",x"c4"),
  2454 => (x"c4",x"1e",x"71",x"31"),
  2455 => (x"92",x"d4",x"4a",x"66"),
  2456 => (x"49",x"c2",x"f8",x"c2"),
  2457 => (x"cd",x"fe",x"81",x"72"),
  2458 => (x"66",x"c4",x"87",x"c5"),
  2459 => (x"e3",x"c0",x"1e",x"49"),
  2460 => (x"dd",x"d6",x"ff",x"49"),
  2461 => (x"ff",x"49",x"d8",x"87"),
  2462 => (x"c8",x"87",x"f2",x"d5"),
  2463 => (x"e6",x"c2",x"1e",x"c0"),
  2464 => (x"e9",x"fd",x"49",x"f2"),
  2465 => (x"d0",x"ff",x"87",x"d5"),
  2466 => (x"78",x"e0",x"c0",x"48"),
  2467 => (x"1e",x"f2",x"e6",x"c2"),
  2468 => (x"d4",x"4a",x"66",x"d0"),
  2469 => (x"c2",x"f8",x"c2",x"92"),
  2470 => (x"fe",x"81",x"72",x"49"),
  2471 => (x"d0",x"87",x"cd",x"cb"),
  2472 => (x"05",x"ac",x"c1",x"86"),
  2473 => (x"c4",x"87",x"cd",x"c1"),
  2474 => (x"31",x"c9",x"49",x"66"),
  2475 => (x"66",x"c4",x"1e",x"71"),
  2476 => (x"c2",x"92",x"d4",x"4a"),
  2477 => (x"72",x"49",x"c2",x"f8"),
  2478 => (x"f2",x"cb",x"fe",x"81"),
  2479 => (x"f2",x"e6",x"c2",x"87"),
  2480 => (x"4a",x"66",x"c8",x"1e"),
  2481 => (x"f8",x"c2",x"92",x"d4"),
  2482 => (x"81",x"72",x"49",x"c2"),
  2483 => (x"87",x"d9",x"c9",x"fe"),
  2484 => (x"1e",x"49",x"66",x"c8"),
  2485 => (x"ff",x"49",x"e3",x"c0"),
  2486 => (x"d7",x"87",x"f7",x"d4"),
  2487 => (x"cc",x"d4",x"ff",x"49"),
  2488 => (x"1e",x"c0",x"c8",x"87"),
  2489 => (x"49",x"f2",x"e6",x"c2"),
  2490 => (x"87",x"d9",x"e7",x"fd"),
  2491 => (x"d0",x"ff",x"86",x"d0"),
  2492 => (x"78",x"e0",x"c0",x"48"),
  2493 => (x"d1",x"fc",x"8e",x"f8"),
  2494 => (x"5b",x"5e",x"0e",x"87"),
  2495 => (x"1e",x"0e",x"5d",x"5c"),
  2496 => (x"d4",x"ff",x"4d",x"71"),
  2497 => (x"7e",x"66",x"d4",x"4c"),
  2498 => (x"a8",x"b7",x"c3",x"48"),
  2499 => (x"c0",x"87",x"c5",x"06"),
  2500 => (x"87",x"e2",x"c1",x"48"),
  2501 => (x"d9",x"fe",x"49",x"75"),
  2502 => (x"1e",x"75",x"87",x"e6"),
  2503 => (x"d4",x"4b",x"66",x"c4"),
  2504 => (x"c2",x"f8",x"c2",x"93"),
  2505 => (x"fe",x"49",x"73",x"83"),
  2506 => (x"c8",x"87",x"e2",x"c4"),
  2507 => (x"ff",x"4b",x"6b",x"83"),
  2508 => (x"e1",x"c8",x"48",x"d0"),
  2509 => (x"73",x"7c",x"dd",x"78"),
  2510 => (x"99",x"ff",x"c3",x"49"),
  2511 => (x"49",x"73",x"7c",x"71"),
  2512 => (x"c3",x"29",x"b7",x"c8"),
  2513 => (x"7c",x"71",x"99",x"ff"),
  2514 => (x"b7",x"d0",x"49",x"73"),
  2515 => (x"99",x"ff",x"c3",x"29"),
  2516 => (x"49",x"73",x"7c",x"71"),
  2517 => (x"71",x"29",x"b7",x"d8"),
  2518 => (x"7c",x"7c",x"c0",x"7c"),
  2519 => (x"7c",x"7c",x"7c",x"7c"),
  2520 => (x"7c",x"7c",x"7c",x"7c"),
  2521 => (x"e0",x"c0",x"7c",x"7c"),
  2522 => (x"1e",x"66",x"c4",x"78"),
  2523 => (x"d2",x"ff",x"49",x"dc"),
  2524 => (x"86",x"c8",x"87",x"e0"),
  2525 => (x"fa",x"26",x"48",x"73"),
  2526 => (x"5e",x"0e",x"87",x"ce"),
  2527 => (x"0e",x"5d",x"5c",x"5b"),
  2528 => (x"ff",x"7e",x"71",x"1e"),
  2529 => (x"1e",x"6e",x"4b",x"d4"),
  2530 => (x"49",x"ea",x"f8",x"c2"),
  2531 => (x"87",x"fd",x"c2",x"fe"),
  2532 => (x"4d",x"70",x"86",x"c4"),
  2533 => (x"c3",x"c3",x"02",x"9d"),
  2534 => (x"f2",x"f8",x"c2",x"87"),
  2535 => (x"49",x"6e",x"4c",x"bf"),
  2536 => (x"87",x"dc",x"d7",x"fe"),
  2537 => (x"c8",x"48",x"d0",x"ff"),
  2538 => (x"d6",x"c1",x"78",x"c5"),
  2539 => (x"15",x"4a",x"c0",x"7b"),
  2540 => (x"c0",x"82",x"c1",x"7b"),
  2541 => (x"04",x"aa",x"b7",x"e0"),
  2542 => (x"d0",x"ff",x"87",x"f5"),
  2543 => (x"c8",x"78",x"c4",x"48"),
  2544 => (x"d3",x"c1",x"78",x"c5"),
  2545 => (x"c4",x"7b",x"c1",x"7b"),
  2546 => (x"02",x"9c",x"74",x"78"),
  2547 => (x"c2",x"87",x"fc",x"c1"),
  2548 => (x"c8",x"7e",x"f2",x"e6"),
  2549 => (x"c0",x"8c",x"4d",x"c0"),
  2550 => (x"c6",x"03",x"ac",x"b7"),
  2551 => (x"a4",x"c0",x"c8",x"87"),
  2552 => (x"c2",x"4c",x"c0",x"4d"),
  2553 => (x"bf",x"97",x"e3",x"f3"),
  2554 => (x"02",x"99",x"d0",x"49"),
  2555 => (x"1e",x"c0",x"87",x"d2"),
  2556 => (x"49",x"ea",x"f8",x"c2"),
  2557 => (x"87",x"f1",x"c4",x"fe"),
  2558 => (x"49",x"70",x"86",x"c4"),
  2559 => (x"87",x"ef",x"c0",x"4a"),
  2560 => (x"1e",x"f2",x"e6",x"c2"),
  2561 => (x"49",x"ea",x"f8",x"c2"),
  2562 => (x"87",x"dd",x"c4",x"fe"),
  2563 => (x"49",x"70",x"86",x"c4"),
  2564 => (x"48",x"d0",x"ff",x"4a"),
  2565 => (x"c1",x"78",x"c5",x"c8"),
  2566 => (x"97",x"6e",x"7b",x"d4"),
  2567 => (x"48",x"6e",x"7b",x"bf"),
  2568 => (x"7e",x"70",x"80",x"c1"),
  2569 => (x"ff",x"05",x"8d",x"c1"),
  2570 => (x"d0",x"ff",x"87",x"f0"),
  2571 => (x"72",x"78",x"c4",x"48"),
  2572 => (x"87",x"c5",x"05",x"9a"),
  2573 => (x"e5",x"c0",x"48",x"c0"),
  2574 => (x"c2",x"1e",x"c1",x"87"),
  2575 => (x"fe",x"49",x"ea",x"f8"),
  2576 => (x"c4",x"87",x"c5",x"c2"),
  2577 => (x"05",x"9c",x"74",x"86"),
  2578 => (x"ff",x"87",x"c4",x"fe"),
  2579 => (x"c5",x"c8",x"48",x"d0"),
  2580 => (x"7b",x"d3",x"c1",x"78"),
  2581 => (x"78",x"c4",x"7b",x"c0"),
  2582 => (x"87",x"c2",x"48",x"c1"),
  2583 => (x"26",x"26",x"48",x"c0"),
  2584 => (x"26",x"4c",x"26",x"4d"),
  2585 => (x"0e",x"4f",x"26",x"4b"),
  2586 => (x"0e",x"5c",x"5b",x"5e"),
  2587 => (x"66",x"cc",x"4b",x"71"),
  2588 => (x"87",x"e7",x"c0",x"02"),
  2589 => (x"8c",x"f0",x"c0",x"4c"),
  2590 => (x"87",x"e6",x"c0",x"02"),
  2591 => (x"8a",x"c1",x"4a",x"74"),
  2592 => (x"8a",x"87",x"df",x"02"),
  2593 => (x"8a",x"87",x"db",x"02"),
  2594 => (x"c0",x"87",x"d7",x"02"),
  2595 => (x"c0",x"02",x"8a",x"e0"),
  2596 => (x"8a",x"c1",x"87",x"e2"),
  2597 => (x"87",x"e3",x"c0",x"02"),
  2598 => (x"73",x"87",x"e5",x"c0"),
  2599 => (x"87",x"da",x"fb",x"49"),
  2600 => (x"1e",x"74",x"87",x"de"),
  2601 => (x"d0",x"f9",x"49",x"c0"),
  2602 => (x"73",x"1e",x"74",x"87"),
  2603 => (x"87",x"c9",x"f9",x"49"),
  2604 => (x"87",x"cc",x"86",x"c8"),
  2605 => (x"e5",x"c1",x"49",x"73"),
  2606 => (x"73",x"87",x"c5",x"87"),
  2607 => (x"87",x"d1",x"c2",x"49"),
  2608 => (x"00",x"87",x"de",x"fe"),
  2609 => (x"c6",x"e6",x"c2",x"1e"),
  2610 => (x"b9",x"c1",x"49",x"bf"),
  2611 => (x"59",x"ca",x"e6",x"c2"),
  2612 => (x"c3",x"48",x"d4",x"ff"),
  2613 => (x"d0",x"ff",x"78",x"ff"),
  2614 => (x"78",x"e1",x"c8",x"48"),
  2615 => (x"c1",x"48",x"d4",x"ff"),
  2616 => (x"71",x"31",x"c4",x"78"),
  2617 => (x"48",x"d0",x"ff",x"78"),
  2618 => (x"26",x"78",x"e0",x"c0"),
  2619 => (x"4a",x"71",x"1e",x"4f"),
  2620 => (x"c2",x"49",x"a2",x"c4"),
  2621 => (x"6a",x"48",x"d9",x"f7"),
  2622 => (x"c1",x"49",x"69",x"78"),
  2623 => (x"ca",x"e6",x"c2",x"b9"),
  2624 => (x"87",x"c0",x"ff",x"59"),
  2625 => (x"87",x"f8",x"cc",x"ff"),
  2626 => (x"4f",x"26",x"48",x"c1"),
  2627 => (x"c4",x"4a",x"71",x"1e"),
  2628 => (x"f7",x"c2",x"49",x"a2"),
  2629 => (x"c2",x"7a",x"bf",x"d9"),
  2630 => (x"79",x"bf",x"c6",x"e6"),
  2631 => (x"71",x"1e",x"4f",x"26"),
  2632 => (x"f8",x"c2",x"1e",x"4a"),
  2633 => (x"fc",x"fd",x"49",x"ea"),
  2634 => (x"86",x"c4",x"87",x"e3"),
  2635 => (x"dc",x"02",x"98",x"70"),
  2636 => (x"f2",x"e6",x"c2",x"87"),
  2637 => (x"ea",x"f8",x"c2",x"1e"),
  2638 => (x"ec",x"ff",x"fd",x"49"),
  2639 => (x"70",x"86",x"c4",x"87"),
  2640 => (x"87",x"c9",x"02",x"98"),
  2641 => (x"49",x"f2",x"e6",x"c2"),
  2642 => (x"c2",x"87",x"e2",x"fe"),
  2643 => (x"26",x"48",x"c0",x"87"),
  2644 => (x"4a",x"71",x"1e",x"4f"),
  2645 => (x"ea",x"f8",x"c2",x"1e"),
  2646 => (x"f0",x"fb",x"fd",x"49"),
  2647 => (x"70",x"86",x"c4",x"87"),
  2648 => (x"87",x"de",x"02",x"98"),
  2649 => (x"49",x"f2",x"e6",x"c2"),
  2650 => (x"c2",x"87",x"e1",x"fe"),
  2651 => (x"c2",x"1e",x"f2",x"e6"),
  2652 => (x"fd",x"49",x"ea",x"f8"),
  2653 => (x"c4",x"87",x"f5",x"ff"),
  2654 => (x"02",x"98",x"70",x"86"),
  2655 => (x"48",x"c1",x"87",x"c4"),
  2656 => (x"48",x"c0",x"87",x"c2"),
  2657 => (x"00",x"00",x"4f",x"26"),
  2658 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

