////////////////////////////////////   MACROS DEFINITIONS  /////////////////////////////////////////
	
`define GUEST_TOP guest_top	// substitute guest_top by guest Mist top module name		

