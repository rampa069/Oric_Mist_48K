library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0f9c287",
    12 => x"86c0c64e",
    13 => x"49c0f9c2",
    14 => x"48cce6c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c7e0",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfcce6",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"e6c21e73",
   176 => x"78c148cc",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"d0e6c287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58d4e6c2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49d4e6",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"e6c287f8",
   280 => x"49bf97d4",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"e6c287e7",
   284 => x"49bf97db",
   285 => x"e6c231d0",
   286 => x"4abf97dc",
   287 => x"b17232c8",
   288 => x"97dde6c2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"dde6c287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97dee6",
   297 => x"2ab7c74a",
   298 => x"e6c2b172",
   299 => x"4abf97d9",
   300 => x"c29dcf4d",
   301 => x"bf97dae6",
   302 => x"ca9ac34a",
   303 => x"dbe6c232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97dce6",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"faeec286",
   323 => x"c278c048",
   324 => x"c01ef2e6",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfcbf2c0",
   331 => x"e8e7c249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f2c07ec0",
   336 => x"c249bfc7",
   337 => x"714ac4e8",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"f8edc287",
   343 => x"eec24dbf",
   344 => x"7ebf9ff0",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bff8edc2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"f2e6c287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f2c087dc",
   358 => x"c249bfc7",
   359 => x"714ac4e8",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"eec287c8",
   363 => x"78c148fa",
   364 => x"f2c087da",
   365 => x"c249bfcb",
   366 => x"714ae8e7",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97f0eec2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"f1eec287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97f2e6",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97fde6",
   387 => x"c0059949",
   388 => x"e6c287cc",
   389 => x"49bf97fe",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97ffe6",
   394 => x"f6eec248",
   395 => x"484c7058",
   396 => x"eec288c1",
   397 => x"e7c258fa",
   398 => x"49bf97c0",
   399 => x"e7c28175",
   400 => x"4abf97c1",
   401 => x"a17232c8",
   402 => x"c7f3c27e",
   403 => x"c2786e48",
   404 => x"bf97c2e7",
   405 => x"58a6c848",
   406 => x"bffaeec2",
   407 => x"87d4c202",
   408 => x"bfc7f2c0",
   409 => x"c4e8c249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"eec287f8",
   415 => x"c24cbff2",
   416 => x"c25cdbf3",
   417 => x"bf97d7e7",
   418 => x"c231c849",
   419 => x"bf97d6e7",
   420 => x"c249a14a",
   421 => x"bf97d8e7",
   422 => x"7232d04a",
   423 => x"e7c249a1",
   424 => x"4abf97d9",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfc7f3c2",
   428 => x"cff3c281",
   429 => x"dfe7c259",
   430 => x"c84abf97",
   431 => x"dee7c232",
   432 => x"a24bbf97",
   433 => x"e0e7c24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97e1e7c2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"d3f3c24a",
   440 => x"cff3c25a",
   441 => x"8ac24abf",
   442 => x"f3c29274",
   443 => x"a17248d3",
   444 => x"87cac178",
   445 => x"97c4e7c2",
   446 => x"31c849bf",
   447 => x"97c3e7c2",
   448 => x"49a14abf",
   449 => x"59c2efc2",
   450 => x"bffeeec2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59dbf3c2",
   454 => x"97c9e7c2",
   455 => x"32c84abf",
   456 => x"97c8e7c2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"d7f3c282",
   460 => x"cff3c25a",
   461 => x"c278c048",
   462 => x"7248cbf3",
   463 => x"f3c278a1",
   464 => x"f3c248db",
   465 => x"c278bfcf",
   466 => x"c248dff3",
   467 => x"78bfd3f3",
   468 => x"bffaeec2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"d7f3c287",
   473 => x"30c448bf",
   474 => x"eec27e70",
   475 => x"786e48fe",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bffaeec2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfc7f3",
   489 => x"bfc3f2c0",
   490 => x"87d902ab",
   491 => x"5bc7f2c0",
   492 => x"1ef2e6c2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"faeec287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81f2e6c2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"e6c291c2",
   505 => x"699f81f2",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"ca49c11e",
   511 => x"86c487ee",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754ac2ef",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c94966c4",
   527 => x"86c487ee",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bffaeec2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48c3f2c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"f6eec2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"eec27b70",
   579 => x"6c49bff2",
   580 => x"757c7181",
   581 => x"f6eec2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"f3c287eb",
   592 => x"c44abfcb",
   593 => x"496949a3",
   594 => x"eec289c2",
   595 => x"7191bff2",
   596 => x"eec24aa2",
   597 => x"6b49bff6",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"cbf3c287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"f2eec289",
   612 => x"a27191bf",
   613 => x"f6eec24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"0e87c9f7",
   620 => x"5d5c5b5e",
   621 => x"4b711e0e",
   622 => x"c94c66d4",
   623 => x"029b732c",
   624 => x"c887cfc1",
   625 => x"026949a3",
   626 => x"d087c7c1",
   627 => x"66d44da3",
   628 => x"f6eec27d",
   629 => x"b9ff49bf",
   630 => x"7e994a6b",
   631 => x"cd03ac71",
   632 => x"7d7bc087",
   633 => x"c44aa3cc",
   634 => x"796a49a3",
   635 => x"8c7287c2",
   636 => x"dd029c74",
   637 => x"731e4987",
   638 => x"87ccfb49",
   639 => x"66d486c4",
   640 => x"99ffc749",
   641 => x"c287cb02",
   642 => x"731ef2e6",
   643 => x"87d9fc49",
   644 => x"f52686c4",
   645 => x"731e87de",
   646 => x"9b4b711e",
   647 => x"87e4c002",
   648 => x"5bdff3c2",
   649 => x"8ac24a73",
   650 => x"bff2eec2",
   651 => x"f3c29249",
   652 => x"7248bfcb",
   653 => x"e3f3c280",
   654 => x"c4487158",
   655 => x"c2efc230",
   656 => x"87edc058",
   657 => x"48dbf3c2",
   658 => x"bfcff3c2",
   659 => x"dff3c278",
   660 => x"d3f3c248",
   661 => x"eec278bf",
   662 => x"c902bffa",
   663 => x"f2eec287",
   664 => x"31c449bf",
   665 => x"f3c287c7",
   666 => x"c449bfd7",
   667 => x"c2efc231",
   668 => x"87c4f459",
   669 => x"5c5b5e0e",
   670 => x"c04a710e",
   671 => x"029a724b",
   672 => x"da87e1c0",
   673 => x"699f49a2",
   674 => x"faeec24b",
   675 => x"87cf02bf",
   676 => x"9f49a2d4",
   677 => x"c04c4969",
   678 => x"d09cffff",
   679 => x"c087c234",
   680 => x"b349744c",
   681 => x"edfd4973",
   682 => x"87caf387",
   683 => x"5c5b5e0e",
   684 => x"86f40e5d",
   685 => x"7ec04a71",
   686 => x"d8029a72",
   687 => x"eee6c287",
   688 => x"c278c048",
   689 => x"c248e6e6",
   690 => x"78bfdff3",
   691 => x"48eae6c2",
   692 => x"bfdbf3c2",
   693 => x"cfefc278",
   694 => x"c250c048",
   695 => x"49bffeee",
   696 => x"bfeee6c2",
   697 => x"03aa714a",
   698 => x"7287ffc3",
   699 => x"0599cf49",
   700 => x"c287e0c0",
   701 => x"c21ef2e6",
   702 => x"49bfe6e6",
   703 => x"48e6e6c2",
   704 => x"7178a1c1",
   705 => x"c487efe3",
   706 => x"fff1c086",
   707 => x"f2e6c248",
   708 => x"c087cc78",
   709 => x"48bffff1",
   710 => x"c080e0c0",
   711 => x"c258c3f2",
   712 => x"48bfeee6",
   713 => x"e6c280c1",
   714 => x"7f2758f2",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e2c202",
   718 => x"02ade5c3",
   719 => x"c087dbc2",
   720 => x"4bbffff1",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181c2ef",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"f9c07ec1",
   744 => x"c8497487",
   745 => x"eac00599",
   746 => x"d0497487",
   747 => x"87d00599",
   748 => x"c00266dc",
   749 => x"497387ca",
   750 => x"700f66dc",
   751 => x"87d30298",
   752 => x"c6c0056e",
   753 => x"c2efc287",
   754 => x"c050c048",
   755 => x"48bffff1",
   756 => x"c287e7c2",
   757 => x"c048cfef",
   758 => x"eec27e50",
   759 => x"c249bffe",
   760 => x"4abfeee6",
   761 => x"fc04aa71",
   762 => x"f3c287c1",
   763 => x"c005bfdf",
   764 => x"eec287c8",
   765 => x"c102bffa",
   766 => x"f2c087fe",
   767 => x"78ff48c3",
   768 => x"bfeae6c2",
   769 => x"87f4ed49",
   770 => x"e6c24970",
   771 => x"a6c459ee",
   772 => x"eae6c248",
   773 => x"eec278bf",
   774 => x"c002bffa",
   775 => x"66c487d8",
   776 => x"ffffcf49",
   777 => x"a999f8ff",
   778 => x"87c5c002",
   779 => x"e1c04dc0",
   780 => x"c04dc187",
   781 => x"66c487dc",
   782 => x"f8ffcf49",
   783 => x"c002a999",
   784 => x"a6c887c8",
   785 => x"c078c048",
   786 => x"a6c887c5",
   787 => x"c878c148",
   788 => x"9d754d66",
   789 => x"87e0c005",
   790 => x"c24966c4",
   791 => x"f2eec289",
   792 => x"c2914abf",
   793 => x"4abfcbf3",
   794 => x"48e6e6c2",
   795 => x"c278a172",
   796 => x"c048eee6",
   797 => x"87e3f978",
   798 => x"8ef448c0",
   799 => x"0087f5eb",
   800 => x"ff000000",
   801 => x"8fffffff",
   802 => x"9800000c",
   803 => x"4600000c",
   804 => x"32335441",
   805 => x"00202020",
   806 => x"31544146",
   807 => x"20202036",
   808 => x"d4ff1e00",
   809 => x"78ffc348",
   810 => x"4f264868",
   811 => x"48d4ff1e",
   812 => x"ff78ffc3",
   813 => x"e1c848d0",
   814 => x"48d4ff78",
   815 => x"f3c278d4",
   816 => x"d4ff48e3",
   817 => x"4f2650bf",
   818 => x"48d0ff1e",
   819 => x"2678e0c0",
   820 => x"ccff1e4f",
   821 => x"99497087",
   822 => x"c087c602",
   823 => x"f105a9fb",
   824 => x"26487187",
   825 => x"5b5e0e4f",
   826 => x"4b710e5c",
   827 => x"f0fe4cc0",
   828 => x"99497087",
   829 => x"87f9c002",
   830 => x"02a9ecc0",
   831 => x"c087f2c0",
   832 => x"c002a9fb",
   833 => x"66cc87eb",
   834 => x"c703acb7",
   835 => x"0266d087",
   836 => x"537187c2",
   837 => x"c2029971",
   838 => x"fe84c187",
   839 => x"497087c3",
   840 => x"87cd0299",
   841 => x"02a9ecc0",
   842 => x"fbc087c7",
   843 => x"d5ff05a9",
   844 => x"0266d087",
   845 => x"97c087c3",
   846 => x"a9ecc07b",
   847 => x"7487c405",
   848 => x"7487c54a",
   849 => x"8a0ac04a",
   850 => x"87c24872",
   851 => x"4c264d26",
   852 => x"4f264b26",
   853 => x"87c9fd1e",
   854 => x"f0c04970",
   855 => x"ca04a9b7",
   856 => x"b7f9c087",
   857 => x"87c301a9",
   858 => x"c189f0c0",
   859 => x"04a9b7c1",
   860 => x"dac187ca",
   861 => x"c301a9b7",
   862 => x"89f7c087",
   863 => x"4f264871",
   864 => x"5c5b5e0e",
   865 => x"ff4a710e",
   866 => x"49724cd4",
   867 => x"7087eac0",
   868 => x"c2029b4b",
   869 => x"ff8bc187",
   870 => x"c5c848d0",
   871 => x"7cd5c178",
   872 => x"31c64973",
   873 => x"97c3e3c2",
   874 => x"71484abf",
   875 => x"ff7c70b0",
   876 => x"78c448d0",
   877 => x"d5fe4873",
   878 => x"5b5e0e87",
   879 => x"f80e5d5c",
   880 => x"c04b7186",
   881 => x"e0fac07e",
   882 => x"df49bf97",
   883 => x"eec005a9",
   884 => x"49a3c887",
   885 => x"c1496997",
   886 => x"dd05a9c3",
   887 => x"49a3c987",
   888 => x"c1496997",
   889 => x"d105a9c6",
   890 => x"49a3ca87",
   891 => x"c1496997",
   892 => x"c505a9c7",
   893 => x"c248c187",
   894 => x"48c087e1",
   895 => x"fa87dcc2",
   896 => x"4cc087ea",
   897 => x"97e0fac0",
   898 => x"a9c049bf",
   899 => x"fa87cf04",
   900 => x"84c187ff",
   901 => x"97e0fac0",
   902 => x"06ac49bf",
   903 => x"fac087f1",
   904 => x"02bf97e0",
   905 => x"f8f987cf",
   906 => x"99497087",
   907 => x"c087c602",
   908 => x"f105a9ec",
   909 => x"f94cc087",
   910 => x"4d7087e7",
   911 => x"c887e2f9",
   912 => x"dcf958a6",
   913 => x"c14a7087",
   914 => x"49a3c884",
   915 => x"ad496997",
   916 => x"c087c702",
   917 => x"c005adff",
   918 => x"a3c987e7",
   919 => x"49699749",
   920 => x"02a966c4",
   921 => x"c04887c7",
   922 => x"d405a8ff",
   923 => x"49a3ca87",
   924 => x"aa496997",
   925 => x"c087c602",
   926 => x"c405aaff",
   927 => x"d07ec187",
   928 => x"adecc087",
   929 => x"c087c602",
   930 => x"c405adfb",
   931 => x"c14cc087",
   932 => x"fe026e7e",
   933 => x"eff887e1",
   934 => x"f8487487",
   935 => x"87ecfa8e",
   936 => x"5b5e0e00",
   937 => x"1e0e5d5c",
   938 => x"4cc04b71",
   939 => x"c004ab4d",
   940 => x"f6c087e8",
   941 => x"9d751ef9",
   942 => x"c087c402",
   943 => x"c187c24a",
   944 => x"ef49724a",
   945 => x"86c487e6",
   946 => x"84c17e70",
   947 => x"87c2056e",
   948 => x"85c14c73",
   949 => x"ff06ac73",
   950 => x"486e87d8",
   951 => x"264d2626",
   952 => x"264b264c",
   953 => x"5b5e0e4f",
   954 => x"1e0e5d5c",
   955 => x"de494c71",
   956 => x"fdf3c291",
   957 => x"9785714d",
   958 => x"ddc1026d",
   959 => x"e8f3c287",
   960 => x"82744abf",
   961 => x"d8fe4972",
   962 => x"6e7e7087",
   963 => x"87f3c002",
   964 => x"4bf0f3c2",
   965 => x"49cb4a6e",
   966 => x"87ccc6ff",
   967 => x"93cb4b74",
   968 => x"83d9e2c1",
   969 => x"fdc083c4",
   970 => x"49747bde",
   971 => x"87d0c7c1",
   972 => x"f3c27b75",
   973 => x"49bf97fc",
   974 => x"f0f3c21e",
   975 => x"e6e4c149",
   976 => x"7486c487",
   977 => x"f7c6c149",
   978 => x"c149c087",
   979 => x"c287d6c8",
   980 => x"c048e4f3",
   981 => x"df49c178",
   982 => x"fd2687fd",
   983 => x"6f4c87ff",
   984 => x"6e696461",
   985 => x"2e2e2e67",
   986 => x"5b5e0e00",
   987 => x"4b710e5c",
   988 => x"e8f3c24a",
   989 => x"497282bf",
   990 => x"7087e6fc",
   991 => x"c4029c4c",
   992 => x"efeb4987",
   993 => x"e8f3c287",
   994 => x"c178c048",
   995 => x"87c7df49",
   996 => x"0e87ccfd",
   997 => x"5d5c5b5e",
   998 => x"c286f40e",
   999 => x"c04df2e6",
  1000 => x"48a6c44c",
  1001 => x"f3c278c0",
  1002 => x"c049bfe8",
  1003 => x"c1c106a9",
  1004 => x"f2e6c287",
  1005 => x"c0029848",
  1006 => x"f6c087f8",
  1007 => x"66c81ef9",
  1008 => x"c487c702",
  1009 => x"78c048a6",
  1010 => x"a6c487c5",
  1011 => x"c478c148",
  1012 => x"d7eb4966",
  1013 => x"7086c487",
  1014 => x"c484c14d",
  1015 => x"80c14866",
  1016 => x"c258a6c8",
  1017 => x"49bfe8f3",
  1018 => x"87c603ac",
  1019 => x"ff059d75",
  1020 => x"4cc087c8",
  1021 => x"c3029d75",
  1022 => x"f6c087e0",
  1023 => x"66c81ef9",
  1024 => x"cc87c702",
  1025 => x"78c048a6",
  1026 => x"a6cc87c5",
  1027 => x"cc78c148",
  1028 => x"d7ea4966",
  1029 => x"7086c487",
  1030 => x"c2026e7e",
  1031 => x"496e87e9",
  1032 => x"699781cb",
  1033 => x"0299d049",
  1034 => x"c087d6c1",
  1035 => x"744ae9fd",
  1036 => x"c191cb49",
  1037 => x"7281d9e2",
  1038 => x"c381c879",
  1039 => x"497451ff",
  1040 => x"f3c291de",
  1041 => x"85714dfd",
  1042 => x"7d97c1c2",
  1043 => x"c049a5c1",
  1044 => x"efc251e0",
  1045 => x"02bf97c2",
  1046 => x"84c187d2",
  1047 => x"c24ba5c2",
  1048 => x"db4ac2ef",
  1049 => x"ffc0ff49",
  1050 => x"87dbc187",
  1051 => x"c049a5cd",
  1052 => x"c284c151",
  1053 => x"4a6e4ba5",
  1054 => x"c0ff49cb",
  1055 => x"c6c187ea",
  1056 => x"e5fbc087",
  1057 => x"cb49744a",
  1058 => x"d9e2c191",
  1059 => x"c2797281",
  1060 => x"bf97c2ef",
  1061 => x"7487d802",
  1062 => x"c191de49",
  1063 => x"fdf3c284",
  1064 => x"c283714b",
  1065 => x"dd4ac2ef",
  1066 => x"fbfffe49",
  1067 => x"7487d887",
  1068 => x"c293de4b",
  1069 => x"cb83fdf3",
  1070 => x"51c049a3",
  1071 => x"6e7384c1",
  1072 => x"fe49cb4a",
  1073 => x"c487e1ff",
  1074 => x"80c14866",
  1075 => x"c758a6c8",
  1076 => x"c5c003ac",
  1077 => x"fc056e87",
  1078 => x"487487e0",
  1079 => x"fcf78ef4",
  1080 => x"1e731e87",
  1081 => x"cb494b71",
  1082 => x"d9e2c191",
  1083 => x"4aa1c881",
  1084 => x"48c3e3c2",
  1085 => x"a1c95012",
  1086 => x"e0fac04a",
  1087 => x"ca501248",
  1088 => x"fcf3c281",
  1089 => x"c2501148",
  1090 => x"bf97fcf3",
  1091 => x"49c01e49",
  1092 => x"87d3ddc1",
  1093 => x"48e4f3c2",
  1094 => x"49c178de",
  1095 => x"2687f8d8",
  1096 => x"1e87fef6",
  1097 => x"cb494a71",
  1098 => x"d9e2c191",
  1099 => x"1181c881",
  1100 => x"e8f3c248",
  1101 => x"e8f3c258",
  1102 => x"c178c048",
  1103 => x"87d7d849",
  1104 => x"c01e4f26",
  1105 => x"dcc0c149",
  1106 => x"1e4f2687",
  1107 => x"d2029971",
  1108 => x"eee3c187",
  1109 => x"f750c048",
  1110 => x"e3c4c180",
  1111 => x"c7e2c140",
  1112 => x"c187ce78",
  1113 => x"c148eae3",
  1114 => x"fc78e8e1",
  1115 => x"c2c5c180",
  1116 => x"0e4f2678",
  1117 => x"0e5c5b5e",
  1118 => x"cb4a4c71",
  1119 => x"d9e2c192",
  1120 => x"49a2c882",
  1121 => x"974ba2c9",
  1122 => x"971e4b6b",
  1123 => x"ca1e4969",
  1124 => x"c0491282",
  1125 => x"c087d7eb",
  1126 => x"87fbd649",
  1127 => x"fdc04974",
  1128 => x"8ef887de",
  1129 => x"1e87f8f4",
  1130 => x"4b711e73",
  1131 => x"87c3ff49",
  1132 => x"fefe4973",
  1133 => x"87e9f487",
  1134 => x"711e731e",
  1135 => x"4aa3c64b",
  1136 => x"c187dc02",
  1137 => x"e4c0028a",
  1138 => x"c1028a87",
  1139 => x"028a87e8",
  1140 => x"8a87cac1",
  1141 => x"87efc002",
  1142 => x"87d9028a",
  1143 => x"c287e9c1",
  1144 => x"df48e4f3",
  1145 => x"d549c178",
  1146 => x"e6c187ed",
  1147 => x"fc49c787",
  1148 => x"dec187f1",
  1149 => x"e8f3c287",
  1150 => x"cbc102bf",
  1151 => x"88c14887",
  1152 => x"58ecf3c2",
  1153 => x"c287c1c1",
  1154 => x"02bfecf3",
  1155 => x"c287f9c0",
  1156 => x"48bfe8f3",
  1157 => x"f3c280c1",
  1158 => x"ebc058ec",
  1159 => x"e8f3c287",
  1160 => x"89c649bf",
  1161 => x"59ecf3c2",
  1162 => x"03a9b7c0",
  1163 => x"f3c287da",
  1164 => x"78c048e8",
  1165 => x"f3c287d2",
  1166 => x"cb02bfec",
  1167 => x"e8f3c287",
  1168 => x"80c648bf",
  1169 => x"58ecf3c2",
  1170 => x"cad449c0",
  1171 => x"c0497387",
  1172 => x"f287edfa",
  1173 => x"5e0e87cb",
  1174 => x"710e5c5b",
  1175 => x"1e66cc4c",
  1176 => x"93cb4b74",
  1177 => x"83d9e2c1",
  1178 => x"6a4aa3c4",
  1179 => x"c7f9fe49",
  1180 => x"e1c3c187",
  1181 => x"49a3c87b",
  1182 => x"c95166d4",
  1183 => x"66d849a3",
  1184 => x"49a3ca51",
  1185 => x"265166dc",
  1186 => x"0e87d4f1",
  1187 => x"5d5c5b5e",
  1188 => x"86d0ff0e",
  1189 => x"c859a6d8",
  1190 => x"78c048a6",
  1191 => x"c4c180fc",
  1192 => x"80c87866",
  1193 => x"80c478c1",
  1194 => x"f3c278c1",
  1195 => x"78c148ec",
  1196 => x"bfe4f3c2",
  1197 => x"de486e7e",
  1198 => x"87cb05a8",
  1199 => x"7087d4f3",
  1200 => x"59a6cc49",
  1201 => x"6e87f8d0",
  1202 => x"05a8df48",
  1203 => x"c187eec1",
  1204 => x"c44966c0",
  1205 => x"c17e6981",
  1206 => x"6e48f4dc",
  1207 => x"4aa1d049",
  1208 => x"aa714120",
  1209 => x"c187f905",
  1210 => x"c14ae1c3",
  1211 => x"7a0a66c0",
  1212 => x"66c0c10a",
  1213 => x"df81c949",
  1214 => x"66c0c151",
  1215 => x"c181ca49",
  1216 => x"c0c151d3",
  1217 => x"81cb4966",
  1218 => x"c44ba1c4",
  1219 => x"786b48a6",
  1220 => x"1e721e71",
  1221 => x"48c4ddc1",
  1222 => x"d04966cc",
  1223 => x"41204aa1",
  1224 => x"f905aa71",
  1225 => x"264a2687",
  1226 => x"c9797249",
  1227 => x"52df4aa1",
  1228 => x"d4c181ca",
  1229 => x"48a6c851",
  1230 => x"c2cf78c2",
  1231 => x"87ece587",
  1232 => x"e587cee6",
  1233 => x"4c7087db",
  1234 => x"02acfbc0",
  1235 => x"d487d0c1",
  1236 => x"c2c10566",
  1237 => x"1e1ec087",
  1238 => x"e4c11ec1",
  1239 => x"49c01ecc",
  1240 => x"c187f3fb",
  1241 => x"c44a66d0",
  1242 => x"c7496a82",
  1243 => x"c1517481",
  1244 => x"6a1ed81e",
  1245 => x"e581c849",
  1246 => x"86d887eb",
  1247 => x"4866c4c1",
  1248 => x"c701a8c0",
  1249 => x"48a6c887",
  1250 => x"87ce78c1",
  1251 => x"4866c4c1",
  1252 => x"a6c888c1",
  1253 => x"e487c358",
  1254 => x"a6cc87f7",
  1255 => x"7478c248",
  1256 => x"d6cd029c",
  1257 => x"4866c887",
  1258 => x"a866c8c1",
  1259 => x"87cbcd03",
  1260 => x"c048a6d8",
  1261 => x"87e9e378",
  1262 => x"d0c14c70",
  1263 => x"d6c205ac",
  1264 => x"7e66d887",
  1265 => x"7087cde6",
  1266 => x"59a6dc49",
  1267 => x"7087d2e3",
  1268 => x"acecc04c",
  1269 => x"87eac105",
  1270 => x"cb4966c8",
  1271 => x"66c0c191",
  1272 => x"4aa1c481",
  1273 => x"a1c84d6a",
  1274 => x"5266d84a",
  1275 => x"79e3c4c1",
  1276 => x"7087eee2",
  1277 => x"d8029c4c",
  1278 => x"acfbc087",
  1279 => x"7487d202",
  1280 => x"87dde255",
  1281 => x"029c4c70",
  1282 => x"fbc087c7",
  1283 => x"eeff05ac",
  1284 => x"55e0c087",
  1285 => x"c055c1c2",
  1286 => x"66d47d97",
  1287 => x"05a96e49",
  1288 => x"66c887db",
  1289 => x"a866c448",
  1290 => x"c887ca04",
  1291 => x"80c14866",
  1292 => x"c858a6cc",
  1293 => x"4866c487",
  1294 => x"a6c888c1",
  1295 => x"87e1e158",
  1296 => x"d0c14c70",
  1297 => x"87c805ac",
  1298 => x"c14866d0",
  1299 => x"58a6d480",
  1300 => x"02acd0c1",
  1301 => x"dc87eafd",
  1302 => x"66d448a6",
  1303 => x"4866d878",
  1304 => x"05a866dc",
  1305 => x"c087e6c9",
  1306 => x"c048a6e0",
  1307 => x"80c478f0",
  1308 => x"c47866cc",
  1309 => x"7e78c080",
  1310 => x"fbc04874",
  1311 => x"a6f0c088",
  1312 => x"02987058",
  1313 => x"4887e1c8",
  1314 => x"f0c088cb",
  1315 => x"987058a6",
  1316 => x"87e9c002",
  1317 => x"c088c948",
  1318 => x"7058a6f0",
  1319 => x"e9c30298",
  1320 => x"88c44887",
  1321 => x"58a6f0c0",
  1322 => x"de029870",
  1323 => x"88c14887",
  1324 => x"58a6f0c0",
  1325 => x"c3029870",
  1326 => x"e5c787d0",
  1327 => x"a6e0c087",
  1328 => x"cc78c048",
  1329 => x"80c14866",
  1330 => x"ff58a6d0",
  1331 => x"7087d2df",
  1332 => x"acecc04c",
  1333 => x"c087d702",
  1334 => x"c00266e0",
  1335 => x"e4c087c7",
  1336 => x"c9c05ca6",
  1337 => x"c0487487",
  1338 => x"e8c088f0",
  1339 => x"ecc058a6",
  1340 => x"cdc002ac",
  1341 => x"e8deff87",
  1342 => x"c04c7087",
  1343 => x"ff05acec",
  1344 => x"e0c087f3",
  1345 => x"66d41e66",
  1346 => x"ecc01e49",
  1347 => x"e4c11e66",
  1348 => x"66d81ecc",
  1349 => x"87fef449",
  1350 => x"1eca1ec0",
  1351 => x"4966e0c0",
  1352 => x"d8c191cb",
  1353 => x"a6d88166",
  1354 => x"78a1c448",
  1355 => x"49bf66d8",
  1356 => x"87f1deff",
  1357 => x"b7c086d8",
  1358 => x"c8c106a8",
  1359 => x"de1ec187",
  1360 => x"bf66c81e",
  1361 => x"dcdeff49",
  1362 => x"7086c887",
  1363 => x"08c04849",
  1364 => x"a6e4c088",
  1365 => x"a8b7c058",
  1366 => x"87e9c006",
  1367 => x"4866e0c0",
  1368 => x"03a8b7dd",
  1369 => x"bf6e87df",
  1370 => x"66e0c049",
  1371 => x"51e0c081",
  1372 => x"81c14966",
  1373 => x"c281bf6e",
  1374 => x"e0c051c1",
  1375 => x"81c24966",
  1376 => x"c081bf6e",
  1377 => x"c47ec151",
  1378 => x"dfff87de",
  1379 => x"e4c087c6",
  1380 => x"deff58a6",
  1381 => x"e8c087fe",
  1382 => x"ecc058a6",
  1383 => x"cbc005a8",
  1384 => x"a6e4c087",
  1385 => x"66e0c048",
  1386 => x"87c4c078",
  1387 => x"87f1dbff",
  1388 => x"cb4966c8",
  1389 => x"66c0c191",
  1390 => x"70807148",
  1391 => x"c84a6e7e",
  1392 => x"ca496e82",
  1393 => x"66e0c081",
  1394 => x"66e4c051",
  1395 => x"c081c149",
  1396 => x"c18966e0",
  1397 => x"70307148",
  1398 => x"7189c149",
  1399 => x"f7c27a97",
  1400 => x"c049bfd9",
  1401 => x"972966e0",
  1402 => x"71484a6a",
  1403 => x"a6f0c098",
  1404 => x"c4496e58",
  1405 => x"dc4d6981",
  1406 => x"66d84866",
  1407 => x"c8c002a8",
  1408 => x"48a6d887",
  1409 => x"c5c078c0",
  1410 => x"48a6d887",
  1411 => x"66d878c1",
  1412 => x"1ee0c01e",
  1413 => x"dbff4975",
  1414 => x"86c887cb",
  1415 => x"b7c04c70",
  1416 => x"d4c106ac",
  1417 => x"c0857487",
  1418 => x"897449e0",
  1419 => x"ddc14b75",
  1420 => x"fe714ad4",
  1421 => x"c287f1e9",
  1422 => x"66e8c085",
  1423 => x"c080c148",
  1424 => x"c058a6ec",
  1425 => x"c14966ec",
  1426 => x"02a97081",
  1427 => x"d887c8c0",
  1428 => x"78c048a6",
  1429 => x"d887c5c0",
  1430 => x"78c148a6",
  1431 => x"c21e66d8",
  1432 => x"e0c049a4",
  1433 => x"70887148",
  1434 => x"49751e49",
  1435 => x"87f5d9ff",
  1436 => x"b7c086c8",
  1437 => x"c0ff01a8",
  1438 => x"66e8c087",
  1439 => x"87d1c002",
  1440 => x"81c9496e",
  1441 => x"5166e8c0",
  1442 => x"c5c1486e",
  1443 => x"ccc078f3",
  1444 => x"c9496e87",
  1445 => x"6e51c281",
  1446 => x"e7c6c148",
  1447 => x"c07ec178",
  1448 => x"d8ff87c6",
  1449 => x"4c7087eb",
  1450 => x"f5c0026e",
  1451 => x"4866c887",
  1452 => x"04a866c4",
  1453 => x"c887cbc0",
  1454 => x"80c14866",
  1455 => x"c058a6cc",
  1456 => x"66c487e0",
  1457 => x"c888c148",
  1458 => x"d5c058a6",
  1459 => x"acc6c187",
  1460 => x"87c8c005",
  1461 => x"c14866cc",
  1462 => x"58a6d080",
  1463 => x"87f1d7ff",
  1464 => x"66d04c70",
  1465 => x"d480c148",
  1466 => x"9c7458a6",
  1467 => x"87cbc002",
  1468 => x"c14866c8",
  1469 => x"04a866c8",
  1470 => x"ff87f5f2",
  1471 => x"c887c9d7",
  1472 => x"a8c74866",
  1473 => x"87e5c003",
  1474 => x"48ecf3c2",
  1475 => x"66c878c0",
  1476 => x"c191cb49",
  1477 => x"c48166c0",
  1478 => x"4a6a4aa1",
  1479 => x"c87952c0",
  1480 => x"80c14866",
  1481 => x"c758a6cc",
  1482 => x"dbff04a8",
  1483 => x"8ed0ff87",
  1484 => x"87e9deff",
  1485 => x"64616f4c",
  1486 => x"74655320",
  1487 => x"676e6974",
  1488 => x"00812073",
  1489 => x"65766153",
  1490 => x"74655320",
  1491 => x"676e6974",
  1492 => x"00812073",
  1493 => x"1e00203a",
  1494 => x"4b711e73",
  1495 => x"87c6029b",
  1496 => x"48e8f3c2",
  1497 => x"1ec778c0",
  1498 => x"bfe8f3c2",
  1499 => x"e2c11e49",
  1500 => x"f3c21ed9",
  1501 => x"ec49bfe4",
  1502 => x"86cc87d1",
  1503 => x"bfe4f3c2",
  1504 => x"87c7e749",
  1505 => x"c8029b73",
  1506 => x"d9e2c187",
  1507 => x"c1e7c049",
  1508 => x"ccddff87",
  1509 => x"1e731e87",
  1510 => x"dfc14bc0",
  1511 => x"c5c149c0",
  1512 => x"e3c287fc",
  1513 => x"50c048c3",
  1514 => x"bffce3c1",
  1515 => x"c9ffc049",
  1516 => x"05987087",
  1517 => x"dfc187c4",
  1518 => x"48734bcc",
  1519 => x"87e1dcff",
  1520 => x"4349524f",
  1521 => x"20202020",
  1522 => x"00474643",
  1523 => x"204d4f52",
  1524 => x"64616f6c",
  1525 => x"20676e69",
  1526 => x"6c696166",
  1527 => x"1e006465",
  1528 => x"c187c8c8",
  1529 => x"87effd49",
  1530 => x"87cfebfe",
  1531 => x"cd029870",
  1532 => x"ccf4fe87",
  1533 => x"02987087",
  1534 => x"4ac187c4",
  1535 => x"4ac087c2",
  1536 => x"ce059a72",
  1537 => x"c11ec087",
  1538 => x"c049efe0",
  1539 => x"c487f9f3",
  1540 => x"c087fe86",
  1541 => x"fae0c11e",
  1542 => x"ebf3c049",
  1543 => x"fd1ec087",
  1544 => x"497087f3",
  1545 => x"87e0f3c0",
  1546 => x"f887ffc3",
  1547 => x"534f268e",
  1548 => x"61662044",
  1549 => x"64656c69",
  1550 => x"6f42002e",
  1551 => x"6e69746f",
  1552 => x"2e2e2e67",
  1553 => x"e8c01e00",
  1554 => x"f7c087eb",
  1555 => x"87f687c5",
  1556 => x"c21e4f26",
  1557 => x"c048e8f3",
  1558 => x"e4f3c278",
  1559 => x"fd78c048",
  1560 => x"87e187fd",
  1561 => x"4f2648c0",
  1562 => x"20202020",
  1563 => x"20202020",
  1564 => x"20202020",
  1565 => x"69784520",
  1566 => x"20202074",
  1567 => x"20202020",
  1568 => x"20202020",
  1569 => x"80008120",
  1570 => x"20202020",
  1571 => x"20202020",
  1572 => x"20202020",
  1573 => x"6b636142",
  1574 => x"00112300",
  1575 => x"002cfd00",
  1576 => x"00000000",
  1577 => x"00001123",
  1578 => x"00002d1b",
  1579 => x"23000000",
  1580 => x"39000011",
  1581 => x"0000002d",
  1582 => x"11230000",
  1583 => x"2d570000",
  1584 => x"00000000",
  1585 => x"00112300",
  1586 => x"002d7500",
  1587 => x"00000000",
  1588 => x"00001123",
  1589 => x"00002d93",
  1590 => x"23000000",
  1591 => x"b1000011",
  1592 => x"0000002d",
  1593 => x"11230000",
  1594 => x"00000000",
  1595 => x"00000000",
  1596 => x"0011b800",
  1597 => x"00000000",
  1598 => x"00000000",
  1599 => x"00001900",
  1600 => x"4349524f",
  1601 => x"20202020",
  1602 => x"004d4f52",
  1603 => x"64616f4c",
  1604 => x"002e2a20",
  1605 => x"48f0fe1e",
  1606 => x"09cd78c0",
  1607 => x"4f260979",
  1608 => x"f0fe1e1e",
  1609 => x"26487ebf",
  1610 => x"fe1e4f26",
  1611 => x"78c148f0",
  1612 => x"fe1e4f26",
  1613 => x"78c048f0",
  1614 => x"711e4f26",
  1615 => x"5252c04a",
  1616 => x"5e0e4f26",
  1617 => x"0e5d5c5b",
  1618 => x"4d7186f4",
  1619 => x"c17e6d97",
  1620 => x"6c974ca5",
  1621 => x"58a6c848",
  1622 => x"66c4486e",
  1623 => x"87c505a8",
  1624 => x"e6c048ff",
  1625 => x"87caff87",
  1626 => x"9749a5c2",
  1627 => x"a3714b6c",
  1628 => x"4b6b974b",
  1629 => x"6e7e6c97",
  1630 => x"c880c148",
  1631 => x"98c758a6",
  1632 => x"7058a6cc",
  1633 => x"e1fe7c97",
  1634 => x"f4487387",
  1635 => x"264d268e",
  1636 => x"264b264c",
  1637 => x"5b5e0e4f",
  1638 => x"86f40e5c",
  1639 => x"66d84c71",
  1640 => x"9affc34a",
  1641 => x"974ba4c2",
  1642 => x"a173496c",
  1643 => x"97517249",
  1644 => x"486e7e6c",
  1645 => x"a6c880c1",
  1646 => x"cc98c758",
  1647 => x"547058a6",
  1648 => x"caff8ef4",
  1649 => x"fd1e1e87",
  1650 => x"bfe087e8",
  1651 => x"e0c0494a",
  1652 => x"cb0299c0",
  1653 => x"c21e7287",
  1654 => x"fe49cff7",
  1655 => x"86c487f7",
  1656 => x"7087fdfc",
  1657 => x"87c2fd7e",
  1658 => x"1e4f2626",
  1659 => x"49cff7c2",
  1660 => x"c187c7fd",
  1661 => x"fc49c5e7",
  1662 => x"d9c587da",
  1663 => x"0e4f2687",
  1664 => x"5d5c5b5e",
  1665 => x"eef7c20e",
  1666 => x"e9c14abf",
  1667 => x"4c49bfd3",
  1668 => x"4d71bc72",
  1669 => x"c087dbfc",
  1670 => x"d049744b",
  1671 => x"87d50299",
  1672 => x"99d04975",
  1673 => x"1ec01e71",
  1674 => x"4ae5efc1",
  1675 => x"49128273",
  1676 => x"c887e4c0",
  1677 => x"2d2cc186",
  1678 => x"04abc883",
  1679 => x"fb87daff",
  1680 => x"e9c187e8",
  1681 => x"f7c248d3",
  1682 => x"2678bfee",
  1683 => x"264c264d",
  1684 => x"004f264b",
  1685 => x"1e000000",
  1686 => x"c848d0ff",
  1687 => x"d4ff78e1",
  1688 => x"c478c548",
  1689 => x"87c30266",
  1690 => x"c878e0c3",
  1691 => x"87c60266",
  1692 => x"c348d4ff",
  1693 => x"d4ff78f0",
  1694 => x"ff787148",
  1695 => x"e1c848d0",
  1696 => x"78e0c078",
  1697 => x"5e0e4f26",
  1698 => x"710e5c5b",
  1699 => x"cff7c24c",
  1700 => x"87eefa49",
  1701 => x"b7c04a70",
  1702 => x"e3c204aa",
  1703 => x"aae0c387",
  1704 => x"c187c905",
  1705 => x"c148c9ed",
  1706 => x"87d4c278",
  1707 => x"05aaf0c3",
  1708 => x"edc187c9",
  1709 => x"78c148c5",
  1710 => x"c187f5c1",
  1711 => x"02bfc9ed",
  1712 => x"4b7287c7",
  1713 => x"c2b3c0c2",
  1714 => x"744b7287",
  1715 => x"87d1059c",
  1716 => x"bfc5edc1",
  1717 => x"c9edc11e",
  1718 => x"49721ebf",
  1719 => x"c887f8fd",
  1720 => x"c5edc186",
  1721 => x"e0c002bf",
  1722 => x"c4497387",
  1723 => x"c19129b7",
  1724 => x"7381e5ee",
  1725 => x"c29acf4a",
  1726 => x"7248c192",
  1727 => x"ff4a7030",
  1728 => x"694872ba",
  1729 => x"db797098",
  1730 => x"c4497387",
  1731 => x"c19129b7",
  1732 => x"7381e5ee",
  1733 => x"c29acf4a",
  1734 => x"7248c392",
  1735 => x"484a7030",
  1736 => x"7970b069",
  1737 => x"48c9edc1",
  1738 => x"edc178c0",
  1739 => x"78c048c5",
  1740 => x"49cff7c2",
  1741 => x"7087cbf8",
  1742 => x"aab7c04a",
  1743 => x"87ddfd03",
  1744 => x"c8fc48c0",
  1745 => x"00000087",
  1746 => x"00000000",
  1747 => x"4a711e00",
  1748 => x"87f2fc49",
  1749 => x"c01e4f26",
  1750 => x"c449724a",
  1751 => x"e5eec191",
  1752 => x"c179c081",
  1753 => x"aab7d082",
  1754 => x"2687ee04",
  1755 => x"5b5e0e4f",
  1756 => x"710e5d5c",
  1757 => x"87faf64d",
  1758 => x"b7c44a75",
  1759 => x"eec1922a",
  1760 => x"4c7582e5",
  1761 => x"94c29ccf",
  1762 => x"744b496a",
  1763 => x"c29bc32b",
  1764 => x"70307448",
  1765 => x"74bcff4c",
  1766 => x"70987148",
  1767 => x"87caf67a",
  1768 => x"e6fa4873",
  1769 => x"00000087",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"261e1600",
  1786 => x"3d362e25",
  1787 => x"d0ff1e3e",
  1788 => x"78e1c848",
  1789 => x"d4ff4871",
  1790 => x"4f267808",
  1791 => x"48d0ff1e",
  1792 => x"7178e1c8",
  1793 => x"08d4ff48",
  1794 => x"4866c478",
  1795 => x"7808d4ff",
  1796 => x"711e4f26",
  1797 => x"4966c44a",
  1798 => x"ff49721e",
  1799 => x"d0ff87de",
  1800 => x"78e0c048",
  1801 => x"1e4f2626",
  1802 => x"b7c24a71",
  1803 => x"87c303aa",
  1804 => x"ce87c282",
  1805 => x"1e66c482",
  1806 => x"d5ff4972",
  1807 => x"4f262687",
  1808 => x"4ad4ff1e",
  1809 => x"ff7affc3",
  1810 => x"e1c848d0",
  1811 => x"c27ade78",
  1812 => x"7abfd9f7",
  1813 => x"28c84849",
  1814 => x"48717a70",
  1815 => x"7a7028d0",
  1816 => x"28d84871",
  1817 => x"d0ff7a70",
  1818 => x"78e0c048",
  1819 => x"5e0e4f26",
  1820 => x"0e5d5c5b",
  1821 => x"f7c24c71",
  1822 => x"4b4dbfd9",
  1823 => x"66d02b74",
  1824 => x"d483c19b",
  1825 => x"c204ab66",
  1826 => x"744bc087",
  1827 => x"4966d04a",
  1828 => x"b9ff3172",
  1829 => x"48739975",
  1830 => x"4a703072",
  1831 => x"c2b07148",
  1832 => x"fe58ddf7",
  1833 => x"4d2687da",
  1834 => x"4b264c26",
  1835 => x"ff1e4f26",
  1836 => x"c9c848d0",
  1837 => x"ff487178",
  1838 => x"267808d4",
  1839 => x"4a711e4f",
  1840 => x"ff87eb49",
  1841 => x"78c848d0",
  1842 => x"731e4f26",
  1843 => x"c24b711e",
  1844 => x"02bfe9f7",
  1845 => x"ebc287c3",
  1846 => x"48d0ff87",
  1847 => x"7378c9c8",
  1848 => x"b1e0c049",
  1849 => x"7148d4ff",
  1850 => x"ddf7c278",
  1851 => x"c878c048",
  1852 => x"87c50266",
  1853 => x"c249ffc3",
  1854 => x"c249c087",
  1855 => x"cc59e5f7",
  1856 => x"87c60266",
  1857 => x"4ad5d5c5",
  1858 => x"ffcf87c4",
  1859 => x"f7c24aff",
  1860 => x"f7c25ae9",
  1861 => x"78c148e9",
  1862 => x"4d2687c4",
  1863 => x"4b264c26",
  1864 => x"5e0e4f26",
  1865 => x"0e5d5c5b",
  1866 => x"f7c24a71",
  1867 => x"724cbfe5",
  1868 => x"87cb029a",
  1869 => x"c191c849",
  1870 => x"714bc0f3",
  1871 => x"c187c483",
  1872 => x"c04bc0f7",
  1873 => x"7449134d",
  1874 => x"e1f7c299",
  1875 => x"d4ffb9bf",
  1876 => x"c1787148",
  1877 => x"c8852cb7",
  1878 => x"e804adb7",
  1879 => x"ddf7c287",
  1880 => x"80c848bf",
  1881 => x"58e1f7c2",
  1882 => x"1e87effe",
  1883 => x"4b711e73",
  1884 => x"029a4a13",
  1885 => x"497287cb",
  1886 => x"1387e7fe",
  1887 => x"f5059a4a",
  1888 => x"87dafe87",
  1889 => x"ddf7c21e",
  1890 => x"f7c249bf",
  1891 => x"a1c148dd",
  1892 => x"b7c0c478",
  1893 => x"87db03a9",
  1894 => x"c248d4ff",
  1895 => x"78bfe1f7",
  1896 => x"bfddf7c2",
  1897 => x"ddf7c249",
  1898 => x"78a1c148",
  1899 => x"a9b7c0c4",
  1900 => x"ff87e504",
  1901 => x"78c848d0",
  1902 => x"48e9f7c2",
  1903 => x"4f2678c0",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"5f000000",
  1907 => x"0000005f",
  1908 => x"00030300",
  1909 => x"00000303",
  1910 => x"147f7f14",
  1911 => x"00147f7f",
  1912 => x"6b2e2400",
  1913 => x"00123a6b",
  1914 => x"18366a4c",
  1915 => x"0032566c",
  1916 => x"594f7e30",
  1917 => x"40683a77",
  1918 => x"07040000",
  1919 => x"00000003",
  1920 => x"3e1c0000",
  1921 => x"00004163",
  1922 => x"63410000",
  1923 => x"00001c3e",
  1924 => x"1c3e2a08",
  1925 => x"082a3e1c",
  1926 => x"3e080800",
  1927 => x"0008083e",
  1928 => x"e0800000",
  1929 => x"00000060",
  1930 => x"08080800",
  1931 => x"00080808",
  1932 => x"60000000",
  1933 => x"00000060",
  1934 => x"18306040",
  1935 => x"0103060c",
  1936 => x"597f3e00",
  1937 => x"003e7f4d",
  1938 => x"7f060400",
  1939 => x"0000007f",
  1940 => x"71634200",
  1941 => x"00464f59",
  1942 => x"49632200",
  1943 => x"00367f49",
  1944 => x"13161c18",
  1945 => x"00107f7f",
  1946 => x"45672700",
  1947 => x"00397d45",
  1948 => x"4b7e3c00",
  1949 => x"00307949",
  1950 => x"71010100",
  1951 => x"00070f79",
  1952 => x"497f3600",
  1953 => x"00367f49",
  1954 => x"494f0600",
  1955 => x"001e3f69",
  1956 => x"66000000",
  1957 => x"00000066",
  1958 => x"e6800000",
  1959 => x"00000066",
  1960 => x"14080800",
  1961 => x"00222214",
  1962 => x"14141400",
  1963 => x"00141414",
  1964 => x"14222200",
  1965 => x"00080814",
  1966 => x"51030200",
  1967 => x"00060f59",
  1968 => x"5d417f3e",
  1969 => x"001e1f55",
  1970 => x"097f7e00",
  1971 => x"007e7f09",
  1972 => x"497f7f00",
  1973 => x"00367f49",
  1974 => x"633e1c00",
  1975 => x"00414141",
  1976 => x"417f7f00",
  1977 => x"001c3e63",
  1978 => x"497f7f00",
  1979 => x"00414149",
  1980 => x"097f7f00",
  1981 => x"00010109",
  1982 => x"417f3e00",
  1983 => x"007a7b49",
  1984 => x"087f7f00",
  1985 => x"007f7f08",
  1986 => x"7f410000",
  1987 => x"0000417f",
  1988 => x"40602000",
  1989 => x"003f7f40",
  1990 => x"1c087f7f",
  1991 => x"00416336",
  1992 => x"407f7f00",
  1993 => x"00404040",
  1994 => x"0c067f7f",
  1995 => x"007f7f06",
  1996 => x"0c067f7f",
  1997 => x"007f7f18",
  1998 => x"417f3e00",
  1999 => x"003e7f41",
  2000 => x"097f7f00",
  2001 => x"00060f09",
  2002 => x"61417f3e",
  2003 => x"00407e7f",
  2004 => x"097f7f00",
  2005 => x"00667f19",
  2006 => x"4d6f2600",
  2007 => x"00327b59",
  2008 => x"7f010100",
  2009 => x"0001017f",
  2010 => x"407f3f00",
  2011 => x"003f7f40",
  2012 => x"703f0f00",
  2013 => x"000f3f70",
  2014 => x"18307f7f",
  2015 => x"007f7f30",
  2016 => x"1c366341",
  2017 => x"4163361c",
  2018 => x"7c060301",
  2019 => x"0103067c",
  2020 => x"4d597161",
  2021 => x"00414347",
  2022 => x"7f7f0000",
  2023 => x"00004141",
  2024 => x"0c060301",
  2025 => x"40603018",
  2026 => x"41410000",
  2027 => x"00007f7f",
  2028 => x"03060c08",
  2029 => x"00080c06",
  2030 => x"80808080",
  2031 => x"00808080",
  2032 => x"03000000",
  2033 => x"00000407",
  2034 => x"54742000",
  2035 => x"00787c54",
  2036 => x"447f7f00",
  2037 => x"00387c44",
  2038 => x"447c3800",
  2039 => x"00004444",
  2040 => x"447c3800",
  2041 => x"007f7f44",
  2042 => x"547c3800",
  2043 => x"00185c54",
  2044 => x"7f7e0400",
  2045 => x"00000505",
  2046 => x"a4bc1800",
  2047 => x"007cfca4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
