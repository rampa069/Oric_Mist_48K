
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"7f",x"7f",x"00"),
     1 => (x"00",x"78",x"7c",x"04"),
     2 => (x"3d",x"00",x"00",x"00"),
     3 => (x"00",x"00",x"40",x"7d"),
     4 => (x"80",x"80",x"80",x"00"),
     5 => (x"00",x"00",x"7d",x"fd"),
     6 => (x"10",x"7f",x"7f",x"00"),
     7 => (x"00",x"44",x"6c",x"38"),
     8 => (x"3f",x"00",x"00",x"00"),
     9 => (x"00",x"00",x"40",x"7f"),
    10 => (x"18",x"0c",x"7c",x"7c"),
    11 => (x"00",x"78",x"7c",x"0c"),
    12 => (x"04",x"7c",x"7c",x"00"),
    13 => (x"00",x"78",x"7c",x"04"),
    14 => (x"44",x"7c",x"38",x"00"),
    15 => (x"00",x"38",x"7c",x"44"),
    16 => (x"24",x"fc",x"fc",x"00"),
    17 => (x"00",x"18",x"3c",x"24"),
    18 => (x"24",x"3c",x"18",x"00"),
    19 => (x"00",x"fc",x"fc",x"24"),
    20 => (x"04",x"7c",x"7c",x"00"),
    21 => (x"00",x"08",x"0c",x"04"),
    22 => (x"54",x"5c",x"48",x"00"),
    23 => (x"00",x"20",x"74",x"54"),
    24 => (x"7f",x"3f",x"04",x"00"),
    25 => (x"00",x"00",x"44",x"44"),
    26 => (x"40",x"7c",x"3c",x"00"),
    27 => (x"00",x"7c",x"7c",x"40"),
    28 => (x"60",x"3c",x"1c",x"00"),
    29 => (x"00",x"1c",x"3c",x"60"),
    30 => (x"30",x"60",x"7c",x"3c"),
    31 => (x"00",x"3c",x"7c",x"60"),
    32 => (x"10",x"38",x"6c",x"44"),
    33 => (x"00",x"44",x"6c",x"38"),
    34 => (x"e0",x"bc",x"1c",x"00"),
    35 => (x"00",x"1c",x"3c",x"60"),
    36 => (x"74",x"64",x"44",x"00"),
    37 => (x"00",x"44",x"4c",x"5c"),
    38 => (x"3e",x"08",x"08",x"00"),
    39 => (x"00",x"41",x"41",x"77"),
    40 => (x"7f",x"00",x"00",x"00"),
    41 => (x"00",x"00",x"00",x"7f"),
    42 => (x"77",x"41",x"41",x"00"),
    43 => (x"00",x"08",x"08",x"3e"),
    44 => (x"03",x"01",x"01",x"02"),
    45 => (x"00",x"01",x"02",x"02"),
    46 => (x"7f",x"7f",x"7f",x"7f"),
    47 => (x"00",x"7f",x"7f",x"7f"),
    48 => (x"1c",x"1c",x"08",x"08"),
    49 => (x"7f",x"7f",x"3e",x"3e"),
    50 => (x"3e",x"3e",x"7f",x"7f"),
    51 => (x"08",x"08",x"1c",x"1c"),
    52 => (x"7c",x"18",x"10",x"00"),
    53 => (x"00",x"10",x"18",x"7c"),
    54 => (x"7c",x"30",x"10",x"00"),
    55 => (x"00",x"10",x"30",x"7c"),
    56 => (x"60",x"60",x"30",x"10"),
    57 => (x"00",x"06",x"1e",x"78"),
    58 => (x"18",x"3c",x"66",x"42"),
    59 => (x"00",x"42",x"66",x"3c"),
    60 => (x"c2",x"6a",x"38",x"78"),
    61 => (x"00",x"38",x"6c",x"c6"),
    62 => (x"60",x"00",x"00",x"60"),
    63 => (x"00",x"60",x"00",x"00"),
    64 => (x"5c",x"5b",x"5e",x"0e"),
    65 => (x"71",x"1e",x"0e",x"5d"),
    66 => (x"fa",x"f7",x"c2",x"4c"),
    67 => (x"4b",x"c0",x"4d",x"bf"),
    68 => (x"ab",x"74",x"1e",x"c0"),
    69 => (x"c4",x"87",x"c7",x"02"),
    70 => (x"78",x"c0",x"48",x"a6"),
    71 => (x"a6",x"c4",x"87",x"c5"),
    72 => (x"c4",x"78",x"c1",x"48"),
    73 => (x"49",x"73",x"1e",x"66"),
    74 => (x"c8",x"87",x"df",x"ee"),
    75 => (x"49",x"e0",x"c0",x"86"),
    76 => (x"c4",x"87",x"ef",x"ef"),
    77 => (x"49",x"6a",x"4a",x"a5"),
    78 => (x"f1",x"87",x"f0",x"f0"),
    79 => (x"85",x"cb",x"87",x"c6"),
    80 => (x"b7",x"c8",x"83",x"c1"),
    81 => (x"c7",x"ff",x"04",x"ab"),
    82 => (x"4d",x"26",x"26",x"87"),
    83 => (x"4b",x"26",x"4c",x"26"),
    84 => (x"71",x"1e",x"4f",x"26"),
    85 => (x"fe",x"f7",x"c2",x"4a"),
    86 => (x"fe",x"f7",x"c2",x"5a"),
    87 => (x"49",x"78",x"c7",x"48"),
    88 => (x"26",x"87",x"dd",x"fe"),
    89 => (x"1e",x"73",x"1e",x"4f"),
    90 => (x"b7",x"c0",x"4a",x"71"),
    91 => (x"87",x"d3",x"03",x"aa"),
    92 => (x"bf",x"f2",x"d5",x"c2"),
    93 => (x"c1",x"87",x"c4",x"05"),
    94 => (x"c0",x"87",x"c2",x"4b"),
    95 => (x"f6",x"d5",x"c2",x"4b"),
    96 => (x"c2",x"87",x"c4",x"5b"),
    97 => (x"c2",x"5a",x"f6",x"d5"),
    98 => (x"4a",x"bf",x"f2",x"d5"),
    99 => (x"c0",x"c1",x"9a",x"c1"),
   100 => (x"e8",x"ec",x"49",x"a2"),
   101 => (x"da",x"d5",x"c2",x"87"),
   102 => (x"d5",x"c2",x"49",x"bf"),
   103 => (x"fc",x"b1",x"bf",x"f2"),
   104 => (x"fe",x"78",x"71",x"48"),
   105 => (x"71",x"1e",x"87",x"e8"),
   106 => (x"1e",x"66",x"c4",x"4a"),
   107 => (x"f6",x"e9",x"49",x"72"),
   108 => (x"4f",x"26",x"26",x"87"),
   109 => (x"f2",x"d5",x"c2",x"1e"),
   110 => (x"d0",x"e6",x"49",x"bf"),
   111 => (x"f2",x"f7",x"c2",x"87"),
   112 => (x"78",x"bf",x"e8",x"48"),
   113 => (x"48",x"ee",x"f7",x"c2"),
   114 => (x"c2",x"78",x"bf",x"ec"),
   115 => (x"4a",x"bf",x"f2",x"f7"),
   116 => (x"99",x"ff",x"c3",x"49"),
   117 => (x"72",x"2a",x"b7",x"c8"),
   118 => (x"c2",x"b0",x"71",x"48"),
   119 => (x"26",x"58",x"fa",x"f7"),
   120 => (x"5b",x"5e",x"0e",x"4f"),
   121 => (x"71",x"0e",x"5d",x"5c"),
   122 => (x"87",x"c8",x"ff",x"4b"),
   123 => (x"48",x"ed",x"f7",x"c2"),
   124 => (x"49",x"73",x"50",x"c0"),
   125 => (x"70",x"87",x"f6",x"e5"),
   126 => (x"9c",x"c2",x"4c",x"49"),
   127 => (x"cd",x"49",x"ee",x"cb"),
   128 => (x"49",x"70",x"87",x"f8"),
   129 => (x"ed",x"f7",x"c2",x"4d"),
   130 => (x"c1",x"05",x"bf",x"97"),
   131 => (x"66",x"d0",x"87",x"e2"),
   132 => (x"f6",x"f7",x"c2",x"49"),
   133 => (x"d6",x"05",x"99",x"bf"),
   134 => (x"49",x"66",x"d4",x"87"),
   135 => (x"bf",x"ee",x"f7",x"c2"),
   136 => (x"87",x"cb",x"05",x"99"),
   137 => (x"c4",x"e5",x"49",x"73"),
   138 => (x"02",x"98",x"70",x"87"),
   139 => (x"c1",x"87",x"c1",x"c1"),
   140 => (x"87",x"c0",x"fe",x"4c"),
   141 => (x"cd",x"cd",x"49",x"75"),
   142 => (x"02",x"98",x"70",x"87"),
   143 => (x"f7",x"c2",x"87",x"c6"),
   144 => (x"50",x"c1",x"48",x"ed"),
   145 => (x"97",x"ed",x"f7",x"c2"),
   146 => (x"e3",x"c0",x"05",x"bf"),
   147 => (x"f6",x"f7",x"c2",x"87"),
   148 => (x"66",x"d0",x"49",x"bf"),
   149 => (x"d6",x"ff",x"05",x"99"),
   150 => (x"ee",x"f7",x"c2",x"87"),
   151 => (x"66",x"d4",x"49",x"bf"),
   152 => (x"ca",x"ff",x"05",x"99"),
   153 => (x"e4",x"49",x"73",x"87"),
   154 => (x"98",x"70",x"87",x"c3"),
   155 => (x"87",x"ff",x"fe",x"05"),
   156 => (x"d5",x"fb",x"48",x"74"),
   157 => (x"5b",x"5e",x"0e",x"87"),
   158 => (x"f8",x"0e",x"5d",x"5c"),
   159 => (x"4c",x"4d",x"c0",x"86"),
   160 => (x"c4",x"7e",x"bf",x"ec"),
   161 => (x"f7",x"c2",x"48",x"a6"),
   162 => (x"c0",x"78",x"bf",x"fa"),
   163 => (x"f7",x"c1",x"1e",x"1e"),
   164 => (x"87",x"cd",x"fd",x"49"),
   165 => (x"98",x"70",x"86",x"c8"),
   166 => (x"87",x"f3",x"c0",x"02"),
   167 => (x"bf",x"da",x"d5",x"c2"),
   168 => (x"c1",x"87",x"c4",x"05"),
   169 => (x"c0",x"87",x"c2",x"7e"),
   170 => (x"da",x"d5",x"c2",x"7e"),
   171 => (x"ca",x"78",x"6e",x"48"),
   172 => (x"66",x"c4",x"1e",x"fc"),
   173 => (x"c4",x"87",x"c9",x"02"),
   174 => (x"d3",x"c2",x"48",x"a6"),
   175 => (x"87",x"c7",x"78",x"f1"),
   176 => (x"c2",x"48",x"a6",x"c4"),
   177 => (x"c4",x"78",x"fc",x"d3"),
   178 => (x"fb",x"c8",x"49",x"66"),
   179 => (x"c1",x"86",x"c4",x"87"),
   180 => (x"c7",x"1e",x"c0",x"1e"),
   181 => (x"87",x"c9",x"fc",x"49"),
   182 => (x"98",x"70",x"86",x"c8"),
   183 => (x"ff",x"87",x"cd",x"02"),
   184 => (x"87",x"c1",x"fa",x"49"),
   185 => (x"e2",x"49",x"da",x"c1"),
   186 => (x"4d",x"c1",x"87",x"c3"),
   187 => (x"97",x"ed",x"f7",x"c2"),
   188 => (x"87",x"c3",x"02",x"bf"),
   189 => (x"c2",x"87",x"cd",x"d7"),
   190 => (x"4b",x"bf",x"f2",x"f7"),
   191 => (x"bf",x"f2",x"d5",x"c2"),
   192 => (x"87",x"e1",x"c1",x"05"),
   193 => (x"bf",x"da",x"d5",x"c2"),
   194 => (x"87",x"f0",x"c0",x"02"),
   195 => (x"c8",x"48",x"a6",x"c4"),
   196 => (x"c2",x"78",x"c0",x"c0"),
   197 => (x"6e",x"7e",x"de",x"d5"),
   198 => (x"6e",x"49",x"bf",x"97"),
   199 => (x"70",x"80",x"c1",x"48"),
   200 => (x"c8",x"e1",x"71",x"7e"),
   201 => (x"02",x"98",x"70",x"87"),
   202 => (x"66",x"c4",x"87",x"c3"),
   203 => (x"48",x"66",x"c4",x"b3"),
   204 => (x"c8",x"28",x"b7",x"c1"),
   205 => (x"98",x"70",x"58",x"a6"),
   206 => (x"87",x"db",x"ff",x"05"),
   207 => (x"e0",x"49",x"fd",x"c3"),
   208 => (x"fa",x"c3",x"87",x"eb"),
   209 => (x"87",x"e5",x"e0",x"49"),
   210 => (x"ff",x"c3",x"49",x"73"),
   211 => (x"c0",x"1e",x"71",x"99"),
   212 => (x"87",x"d2",x"f9",x"49"),
   213 => (x"b7",x"c8",x"49",x"73"),
   214 => (x"c1",x"1e",x"71",x"29"),
   215 => (x"87",x"c6",x"f9",x"49"),
   216 => (x"c7",x"c6",x"86",x"c8"),
   217 => (x"f6",x"f7",x"c2",x"87"),
   218 => (x"02",x"9b",x"4b",x"bf"),
   219 => (x"d5",x"c2",x"87",x"df"),
   220 => (x"c8",x"49",x"bf",x"ee"),
   221 => (x"98",x"70",x"87",x"d0"),
   222 => (x"87",x"c4",x"c0",x"05"),
   223 => (x"87",x"d3",x"4b",x"c0"),
   224 => (x"c7",x"49",x"e0",x"c2"),
   225 => (x"d5",x"c2",x"87",x"f4"),
   226 => (x"c6",x"c0",x"58",x"f2"),
   227 => (x"ee",x"d5",x"c2",x"87"),
   228 => (x"73",x"78",x"c0",x"48"),
   229 => (x"05",x"99",x"c2",x"49"),
   230 => (x"c3",x"87",x"cf",x"c0"),
   231 => (x"df",x"ff",x"49",x"eb"),
   232 => (x"49",x"70",x"87",x"cb"),
   233 => (x"c0",x"02",x"99",x"c2"),
   234 => (x"4c",x"fb",x"87",x"c2"),
   235 => (x"99",x"c1",x"49",x"73"),
   236 => (x"87",x"cf",x"c0",x"05"),
   237 => (x"ff",x"49",x"f4",x"c3"),
   238 => (x"70",x"87",x"f2",x"de"),
   239 => (x"02",x"99",x"c2",x"49"),
   240 => (x"fa",x"87",x"c2",x"c0"),
   241 => (x"c8",x"49",x"73",x"4c"),
   242 => (x"cf",x"c0",x"05",x"99"),
   243 => (x"49",x"f5",x"c3",x"87"),
   244 => (x"87",x"d9",x"de",x"ff"),
   245 => (x"99",x"c2",x"49",x"70"),
   246 => (x"87",x"d6",x"c0",x"02"),
   247 => (x"bf",x"fe",x"f7",x"c2"),
   248 => (x"87",x"ca",x"c0",x"02"),
   249 => (x"c2",x"88",x"c1",x"48"),
   250 => (x"c0",x"58",x"c2",x"f8"),
   251 => (x"4c",x"ff",x"87",x"c2"),
   252 => (x"49",x"73",x"4d",x"c1"),
   253 => (x"c0",x"05",x"99",x"c4"),
   254 => (x"f2",x"c3",x"87",x"cf"),
   255 => (x"ec",x"dd",x"ff",x"49"),
   256 => (x"c2",x"49",x"70",x"87"),
   257 => (x"dc",x"c0",x"02",x"99"),
   258 => (x"fe",x"f7",x"c2",x"87"),
   259 => (x"c7",x"48",x"7e",x"bf"),
   260 => (x"c0",x"03",x"a8",x"b7"),
   261 => (x"48",x"6e",x"87",x"cb"),
   262 => (x"f8",x"c2",x"80",x"c1"),
   263 => (x"c2",x"c0",x"58",x"c2"),
   264 => (x"c1",x"4c",x"fe",x"87"),
   265 => (x"49",x"fd",x"c3",x"4d"),
   266 => (x"87",x"c1",x"dd",x"ff"),
   267 => (x"99",x"c2",x"49",x"70"),
   268 => (x"87",x"d5",x"c0",x"02"),
   269 => (x"bf",x"fe",x"f7",x"c2"),
   270 => (x"87",x"c9",x"c0",x"02"),
   271 => (x"48",x"fe",x"f7",x"c2"),
   272 => (x"c2",x"c0",x"78",x"c0"),
   273 => (x"c1",x"4c",x"fd",x"87"),
   274 => (x"49",x"fa",x"c3",x"4d"),
   275 => (x"87",x"dd",x"dc",x"ff"),
   276 => (x"99",x"c2",x"49",x"70"),
   277 => (x"87",x"d9",x"c0",x"02"),
   278 => (x"bf",x"fe",x"f7",x"c2"),
   279 => (x"a8",x"b7",x"c7",x"48"),
   280 => (x"87",x"c9",x"c0",x"03"),
   281 => (x"48",x"fe",x"f7",x"c2"),
   282 => (x"c2",x"c0",x"78",x"c7"),
   283 => (x"c1",x"4c",x"fc",x"87"),
   284 => (x"ac",x"b7",x"c0",x"4d"),
   285 => (x"87",x"d5",x"c0",x"03"),
   286 => (x"c1",x"48",x"66",x"c4"),
   287 => (x"7e",x"70",x"80",x"d8"),
   288 => (x"c0",x"02",x"bf",x"6e"),
   289 => (x"bf",x"6e",x"87",x"c7"),
   290 => (x"73",x"49",x"74",x"4b"),
   291 => (x"c3",x"1e",x"c0",x"0f"),
   292 => (x"da",x"c1",x"1e",x"f0"),
   293 => (x"87",x"c9",x"f5",x"49"),
   294 => (x"98",x"70",x"86",x"c8"),
   295 => (x"87",x"d9",x"c0",x"02"),
   296 => (x"bf",x"fe",x"f7",x"c2"),
   297 => (x"cb",x"49",x"6e",x"7e"),
   298 => (x"4a",x"66",x"c4",x"91"),
   299 => (x"02",x"6a",x"82",x"71"),
   300 => (x"6a",x"87",x"c6",x"c0"),
   301 => (x"73",x"49",x"6e",x"4b"),
   302 => (x"02",x"9d",x"75",x"0f"),
   303 => (x"c2",x"87",x"c8",x"c0"),
   304 => (x"49",x"bf",x"fe",x"f7"),
   305 => (x"c2",x"87",x"f9",x"f0"),
   306 => (x"02",x"bf",x"f6",x"d5"),
   307 => (x"49",x"87",x"dd",x"c0"),
   308 => (x"70",x"87",x"f3",x"c2"),
   309 => (x"d3",x"c0",x"02",x"98"),
   310 => (x"fe",x"f7",x"c2",x"87"),
   311 => (x"df",x"f0",x"49",x"bf"),
   312 => (x"f1",x"49",x"c0",x"87"),
   313 => (x"d5",x"c2",x"87",x"ff"),
   314 => (x"78",x"c0",x"48",x"f6"),
   315 => (x"d9",x"f1",x"8e",x"f8"),
   316 => (x"79",x"6f",x"4a",x"87"),
   317 => (x"73",x"79",x"65",x"6b"),
   318 => (x"00",x"6e",x"6f",x"20"),
   319 => (x"6b",x"79",x"6f",x"4a"),
   320 => (x"20",x"73",x"79",x"65"),
   321 => (x"00",x"66",x"66",x"6f"),
   322 => (x"5c",x"5b",x"5e",x"0e"),
   323 => (x"71",x"1e",x"0e",x"5d"),
   324 => (x"fa",x"f7",x"c2",x"4c"),
   325 => (x"cd",x"c1",x"49",x"bf"),
   326 => (x"d1",x"c1",x"4d",x"a1"),
   327 => (x"74",x"7e",x"69",x"81"),
   328 => (x"87",x"cf",x"02",x"9c"),
   329 => (x"74",x"4b",x"a5",x"c4"),
   330 => (x"fa",x"f7",x"c2",x"7b"),
   331 => (x"e1",x"f0",x"49",x"bf"),
   332 => (x"74",x"7b",x"6e",x"87"),
   333 => (x"87",x"c4",x"05",x"9c"),
   334 => (x"87",x"c2",x"4b",x"c0"),
   335 => (x"49",x"73",x"4b",x"c1"),
   336 => (x"d4",x"87",x"e2",x"f0"),
   337 => (x"87",x"c8",x"02",x"66"),
   338 => (x"87",x"ee",x"c0",x"49"),
   339 => (x"87",x"c2",x"4a",x"70"),
   340 => (x"d5",x"c2",x"4a",x"c0"),
   341 => (x"ef",x"26",x"5a",x"fa"),
   342 => (x"00",x"00",x"87",x"f0"),
   343 => (x"12",x"58",x"00",x"00"),
   344 => (x"1b",x"1d",x"14",x"11"),
   345 => (x"59",x"5a",x"23",x"1c"),
   346 => (x"f2",x"f5",x"94",x"91"),
   347 => (x"00",x"00",x"f4",x"eb"),
   348 => (x"00",x"00",x"00",x"00"),
   349 => (x"00",x"00",x"00",x"00"),
   350 => (x"71",x"1e",x"00",x"00"),
   351 => (x"bf",x"c8",x"ff",x"4a"),
   352 => (x"48",x"a1",x"72",x"49"),
   353 => (x"ff",x"1e",x"4f",x"26"),
   354 => (x"fe",x"89",x"bf",x"c8"),
   355 => (x"c0",x"c0",x"c0",x"c0"),
   356 => (x"c4",x"01",x"a9",x"c0"),
   357 => (x"c2",x"4a",x"c0",x"87"),
   358 => (x"72",x"4a",x"c1",x"87"),
   359 => (x"0e",x"4f",x"26",x"48"),
   360 => (x"5d",x"5c",x"5b",x"5e"),
   361 => (x"ff",x"4b",x"71",x"0e"),
   362 => (x"66",x"d0",x"4c",x"d4"),
   363 => (x"d6",x"78",x"c0",x"48"),
   364 => (x"f8",x"d8",x"ff",x"49"),
   365 => (x"7c",x"ff",x"c3",x"87"),
   366 => (x"ff",x"c3",x"49",x"6c"),
   367 => (x"49",x"4d",x"71",x"99"),
   368 => (x"c1",x"99",x"f0",x"c3"),
   369 => (x"cb",x"05",x"a9",x"e0"),
   370 => (x"7c",x"ff",x"c3",x"87"),
   371 => (x"98",x"c3",x"48",x"6c"),
   372 => (x"78",x"08",x"66",x"d0"),
   373 => (x"6c",x"7c",x"ff",x"c3"),
   374 => (x"31",x"c8",x"49",x"4a"),
   375 => (x"6c",x"7c",x"ff",x"c3"),
   376 => (x"72",x"b2",x"71",x"4a"),
   377 => (x"c3",x"31",x"c8",x"49"),
   378 => (x"4a",x"6c",x"7c",x"ff"),
   379 => (x"49",x"72",x"b2",x"71"),
   380 => (x"ff",x"c3",x"31",x"c8"),
   381 => (x"71",x"4a",x"6c",x"7c"),
   382 => (x"48",x"d0",x"ff",x"b2"),
   383 => (x"73",x"78",x"e0",x"c0"),
   384 => (x"87",x"c2",x"02",x"9b"),
   385 => (x"48",x"75",x"7b",x"72"),
   386 => (x"4c",x"26",x"4d",x"26"),
   387 => (x"4f",x"26",x"4b",x"26"),
   388 => (x"0e",x"4f",x"26",x"1e"),
   389 => (x"0e",x"5c",x"5b",x"5e"),
   390 => (x"1e",x"76",x"86",x"f8"),
   391 => (x"fd",x"49",x"a6",x"c8"),
   392 => (x"86",x"c4",x"87",x"fd"),
   393 => (x"48",x"6e",x"4b",x"70"),
   394 => (x"c3",x"03",x"a8",x"c2"),
   395 => (x"4a",x"73",x"87",x"c6"),
   396 => (x"c1",x"9a",x"f0",x"c3"),
   397 => (x"c7",x"02",x"aa",x"d0"),
   398 => (x"aa",x"e0",x"c1",x"87"),
   399 => (x"87",x"f4",x"c2",x"05"),
   400 => (x"99",x"c8",x"49",x"73"),
   401 => (x"ff",x"87",x"c3",x"02"),
   402 => (x"4c",x"73",x"87",x"c6"),
   403 => (x"ac",x"c2",x"9c",x"c3"),
   404 => (x"87",x"cd",x"c1",x"05"),
   405 => (x"c9",x"49",x"66",x"c4"),
   406 => (x"c4",x"1e",x"71",x"31"),
   407 => (x"92",x"d4",x"4a",x"66"),
   408 => (x"49",x"c2",x"f8",x"c2"),
   409 => (x"cd",x"fe",x"81",x"72"),
   410 => (x"66",x"c4",x"87",x"c5"),
   411 => (x"e3",x"c0",x"1e",x"49"),
   412 => (x"dd",x"d6",x"ff",x"49"),
   413 => (x"ff",x"49",x"d8",x"87"),
   414 => (x"c8",x"87",x"f2",x"d5"),
   415 => (x"e6",x"c2",x"1e",x"c0"),
   416 => (x"e9",x"fd",x"49",x"f2"),
   417 => (x"d0",x"ff",x"87",x"d5"),
   418 => (x"78",x"e0",x"c0",x"48"),
   419 => (x"1e",x"f2",x"e6",x"c2"),
   420 => (x"d4",x"4a",x"66",x"d0"),
   421 => (x"c2",x"f8",x"c2",x"92"),
   422 => (x"fe",x"81",x"72",x"49"),
   423 => (x"d0",x"87",x"cd",x"cb"),
   424 => (x"05",x"ac",x"c1",x"86"),
   425 => (x"c4",x"87",x"cd",x"c1"),
   426 => (x"31",x"c9",x"49",x"66"),
   427 => (x"66",x"c4",x"1e",x"71"),
   428 => (x"c2",x"92",x"d4",x"4a"),
   429 => (x"72",x"49",x"c2",x"f8"),
   430 => (x"f2",x"cb",x"fe",x"81"),
   431 => (x"f2",x"e6",x"c2",x"87"),
   432 => (x"4a",x"66",x"c8",x"1e"),
   433 => (x"f8",x"c2",x"92",x"d4"),
   434 => (x"81",x"72",x"49",x"c2"),
   435 => (x"87",x"d9",x"c9",x"fe"),
   436 => (x"1e",x"49",x"66",x"c8"),
   437 => (x"ff",x"49",x"e3",x"c0"),
   438 => (x"d7",x"87",x"f7",x"d4"),
   439 => (x"cc",x"d4",x"ff",x"49"),
   440 => (x"1e",x"c0",x"c8",x"87"),
   441 => (x"49",x"f2",x"e6",x"c2"),
   442 => (x"87",x"d9",x"e7",x"fd"),
   443 => (x"d0",x"ff",x"86",x"d0"),
   444 => (x"78",x"e0",x"c0",x"48"),
   445 => (x"d1",x"fc",x"8e",x"f8"),
   446 => (x"5b",x"5e",x"0e",x"87"),
   447 => (x"1e",x"0e",x"5d",x"5c"),
   448 => (x"d4",x"ff",x"4d",x"71"),
   449 => (x"7e",x"66",x"d4",x"4c"),
   450 => (x"a8",x"b7",x"c3",x"48"),
   451 => (x"c0",x"87",x"c5",x"06"),
   452 => (x"87",x"e2",x"c1",x"48"),
   453 => (x"d9",x"fe",x"49",x"75"),
   454 => (x"1e",x"75",x"87",x"e6"),
   455 => (x"d4",x"4b",x"66",x"c4"),
   456 => (x"c2",x"f8",x"c2",x"93"),
   457 => (x"fe",x"49",x"73",x"83"),
   458 => (x"c8",x"87",x"e2",x"c4"),
   459 => (x"ff",x"4b",x"6b",x"83"),
   460 => (x"e1",x"c8",x"48",x"d0"),
   461 => (x"73",x"7c",x"dd",x"78"),
   462 => (x"99",x"ff",x"c3",x"49"),
   463 => (x"49",x"73",x"7c",x"71"),
   464 => (x"c3",x"29",x"b7",x"c8"),
   465 => (x"7c",x"71",x"99",x"ff"),
   466 => (x"b7",x"d0",x"49",x"73"),
   467 => (x"99",x"ff",x"c3",x"29"),
   468 => (x"49",x"73",x"7c",x"71"),
   469 => (x"71",x"29",x"b7",x"d8"),
   470 => (x"7c",x"7c",x"c0",x"7c"),
   471 => (x"7c",x"7c",x"7c",x"7c"),
   472 => (x"7c",x"7c",x"7c",x"7c"),
   473 => (x"e0",x"c0",x"7c",x"7c"),
   474 => (x"1e",x"66",x"c4",x"78"),
   475 => (x"d2",x"ff",x"49",x"dc"),
   476 => (x"86",x"c8",x"87",x"e0"),
   477 => (x"fa",x"26",x"48",x"73"),
   478 => (x"5e",x"0e",x"87",x"ce"),
   479 => (x"0e",x"5d",x"5c",x"5b"),
   480 => (x"ff",x"7e",x"71",x"1e"),
   481 => (x"1e",x"6e",x"4b",x"d4"),
   482 => (x"49",x"ea",x"f8",x"c2"),
   483 => (x"87",x"fd",x"c2",x"fe"),
   484 => (x"4d",x"70",x"86",x"c4"),
   485 => (x"c3",x"c3",x"02",x"9d"),
   486 => (x"f2",x"f8",x"c2",x"87"),
   487 => (x"49",x"6e",x"4c",x"bf"),
   488 => (x"87",x"dc",x"d7",x"fe"),
   489 => (x"c8",x"48",x"d0",x"ff"),
   490 => (x"d6",x"c1",x"78",x"c5"),
   491 => (x"15",x"4a",x"c0",x"7b"),
   492 => (x"c0",x"82",x"c1",x"7b"),
   493 => (x"04",x"aa",x"b7",x"e0"),
   494 => (x"d0",x"ff",x"87",x"f5"),
   495 => (x"c8",x"78",x"c4",x"48"),
   496 => (x"d3",x"c1",x"78",x"c5"),
   497 => (x"c4",x"7b",x"c1",x"7b"),
   498 => (x"02",x"9c",x"74",x"78"),
   499 => (x"c2",x"87",x"fc",x"c1"),
   500 => (x"c8",x"7e",x"f2",x"e6"),
   501 => (x"c0",x"8c",x"4d",x"c0"),
   502 => (x"c6",x"03",x"ac",x"b7"),
   503 => (x"a4",x"c0",x"c8",x"87"),
   504 => (x"c2",x"4c",x"c0",x"4d"),
   505 => (x"bf",x"97",x"e3",x"f3"),
   506 => (x"02",x"99",x"d0",x"49"),
   507 => (x"1e",x"c0",x"87",x"d2"),
   508 => (x"49",x"ea",x"f8",x"c2"),
   509 => (x"87",x"f1",x"c4",x"fe"),
   510 => (x"49",x"70",x"86",x"c4"),
   511 => (x"87",x"ef",x"c0",x"4a"),
   512 => (x"1e",x"f2",x"e6",x"c2"),
   513 => (x"49",x"ea",x"f8",x"c2"),
   514 => (x"87",x"dd",x"c4",x"fe"),
   515 => (x"49",x"70",x"86",x"c4"),
   516 => (x"48",x"d0",x"ff",x"4a"),
   517 => (x"c1",x"78",x"c5",x"c8"),
   518 => (x"97",x"6e",x"7b",x"d4"),
   519 => (x"48",x"6e",x"7b",x"bf"),
   520 => (x"7e",x"70",x"80",x"c1"),
   521 => (x"ff",x"05",x"8d",x"c1"),
   522 => (x"d0",x"ff",x"87",x"f0"),
   523 => (x"72",x"78",x"c4",x"48"),
   524 => (x"87",x"c5",x"05",x"9a"),
   525 => (x"e5",x"c0",x"48",x"c0"),
   526 => (x"c2",x"1e",x"c1",x"87"),
   527 => (x"fe",x"49",x"ea",x"f8"),
   528 => (x"c4",x"87",x"c5",x"c2"),
   529 => (x"05",x"9c",x"74",x"86"),
   530 => (x"ff",x"87",x"c4",x"fe"),
   531 => (x"c5",x"c8",x"48",x"d0"),
   532 => (x"7b",x"d3",x"c1",x"78"),
   533 => (x"78",x"c4",x"7b",x"c0"),
   534 => (x"87",x"c2",x"48",x"c1"),
   535 => (x"26",x"26",x"48",x"c0"),
   536 => (x"26",x"4c",x"26",x"4d"),
   537 => (x"0e",x"4f",x"26",x"4b"),
   538 => (x"0e",x"5c",x"5b",x"5e"),
   539 => (x"66",x"cc",x"4b",x"71"),
   540 => (x"87",x"e7",x"c0",x"02"),
   541 => (x"8c",x"f0",x"c0",x"4c"),
   542 => (x"87",x"e6",x"c0",x"02"),
   543 => (x"8a",x"c1",x"4a",x"74"),
   544 => (x"8a",x"87",x"df",x"02"),
   545 => (x"8a",x"87",x"db",x"02"),
   546 => (x"c0",x"87",x"d7",x"02"),
   547 => (x"c0",x"02",x"8a",x"e0"),
   548 => (x"8a",x"c1",x"87",x"e2"),
   549 => (x"87",x"e3",x"c0",x"02"),
   550 => (x"73",x"87",x"e5",x"c0"),
   551 => (x"87",x"da",x"fb",x"49"),
   552 => (x"1e",x"74",x"87",x"de"),
   553 => (x"d0",x"f9",x"49",x"c0"),
   554 => (x"73",x"1e",x"74",x"87"),
   555 => (x"87",x"c9",x"f9",x"49"),
   556 => (x"87",x"cc",x"86",x"c8"),
   557 => (x"e5",x"c1",x"49",x"73"),
   558 => (x"73",x"87",x"c5",x"87"),
   559 => (x"87",x"d1",x"c2",x"49"),
   560 => (x"00",x"87",x"de",x"fe"),
   561 => (x"c6",x"e6",x"c2",x"1e"),
   562 => (x"b9",x"c1",x"49",x"bf"),
   563 => (x"59",x"ca",x"e6",x"c2"),
   564 => (x"c3",x"48",x"d4",x"ff"),
   565 => (x"d0",x"ff",x"78",x"ff"),
   566 => (x"78",x"e1",x"c8",x"48"),
   567 => (x"c1",x"48",x"d4",x"ff"),
   568 => (x"71",x"31",x"c4",x"78"),
   569 => (x"48",x"d0",x"ff",x"78"),
   570 => (x"26",x"78",x"e0",x"c0"),
   571 => (x"4a",x"71",x"1e",x"4f"),
   572 => (x"c2",x"49",x"a2",x"c4"),
   573 => (x"6a",x"48",x"d9",x"f7"),
   574 => (x"c1",x"49",x"69",x"78"),
   575 => (x"ca",x"e6",x"c2",x"b9"),
   576 => (x"87",x"c0",x"ff",x"59"),
   577 => (x"87",x"f8",x"cc",x"ff"),
   578 => (x"4f",x"26",x"48",x"c1"),
   579 => (x"c4",x"4a",x"71",x"1e"),
   580 => (x"f7",x"c2",x"49",x"a2"),
   581 => (x"c2",x"7a",x"bf",x"d9"),
   582 => (x"79",x"bf",x"c6",x"e6"),
   583 => (x"71",x"1e",x"4f",x"26"),
   584 => (x"f8",x"c2",x"1e",x"4a"),
   585 => (x"fc",x"fd",x"49",x"ea"),
   586 => (x"86",x"c4",x"87",x"e3"),
   587 => (x"dc",x"02",x"98",x"70"),
   588 => (x"f2",x"e6",x"c2",x"87"),
   589 => (x"ea",x"f8",x"c2",x"1e"),
   590 => (x"ec",x"ff",x"fd",x"49"),
   591 => (x"70",x"86",x"c4",x"87"),
   592 => (x"87",x"c9",x"02",x"98"),
   593 => (x"49",x"f2",x"e6",x"c2"),
   594 => (x"c2",x"87",x"e2",x"fe"),
   595 => (x"26",x"48",x"c0",x"87"),
   596 => (x"4a",x"71",x"1e",x"4f"),
   597 => (x"ea",x"f8",x"c2",x"1e"),
   598 => (x"f0",x"fb",x"fd",x"49"),
   599 => (x"70",x"86",x"c4",x"87"),
   600 => (x"87",x"de",x"02",x"98"),
   601 => (x"49",x"f2",x"e6",x"c2"),
   602 => (x"c2",x"87",x"e1",x"fe"),
   603 => (x"c2",x"1e",x"f2",x"e6"),
   604 => (x"fd",x"49",x"ea",x"f8"),
   605 => (x"c4",x"87",x"f5",x"ff"),
   606 => (x"02",x"98",x"70",x"86"),
   607 => (x"48",x"c1",x"87",x"c4"),
   608 => (x"48",x"c0",x"87",x"c2"),
   609 => (x"00",x"00",x"4f",x"26"),
   610 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

