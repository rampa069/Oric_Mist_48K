--
-- Multicore 2 / Multicore 2+
--
-- Copyright (c) 2017-2020 - Victor Trucco
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS CODE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- You are responsible for any legal issues arising from your use of this code.
--
		
library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity vga_font is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic
);
end entity;

architecture prom of vga_font is
	type rom is array(0 to  16383) of std_logic;
	signal rom_data: rom := (
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','1','1','0','1','0','0','0','0','0','0','0','1','0',
		'1','0','0','0','0','0','0','0','1','0','0','0','0','0','1','0',
		'0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0',
		'1','0','0','0','0','0','1','0','0','0','0','0','0','0','1','0',
		'1','0','0','0','0','0','0','0','1','0','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','1','1','0','0','1','1','1','1','1','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','1','1','0','0','1','1','1','1','1','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','1','0','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','0','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','1','1','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','1','0','1','1','0','1','1','0','1','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1',
		'0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','1','1','1','1','1','1','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','0','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0',
		'0','0','1','1','1','1','0','0','0','1','1','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','1','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','1','1','1','1','0','1','1','0','1','1','1','1','0',
		'1','1','0','1','1','1','1','0','1','1','0','1','1','1','0','0',
		'1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','1','0',
		'0','1','1','0','0','1','1','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','1','1','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','0','1','0','0','1','1','0','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','0','1','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','0','1','0','0','1','1','0','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','0','1','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','1','1','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','0','1','1','1','0','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','1','1','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','0','1','1','1','0',
		'1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'1','1','1','1','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','1','1','1','1','0','1','1','0','0','1','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','1','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0',
		'0','1','0','1','1','0','1','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','0','1','1','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','1','0','1','1','1','0','0','1','1','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','1','1','0',
		'1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0',
		'0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','1','1','1','1','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','0','0','0','1','1','0','0','0','0','0',
		'1','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','0','1','1','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','1','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','1','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','0','1','1','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','1','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','1','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','0','1','1','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','1','1','1','0','0',
		'0','1','1','1','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','1','1','1','1','1','1','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','1','1','0','0','0','0','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','1','1','1','1','1','0','0','1','1','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','0','1','1','1','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0',
		'1','1','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','0','1','1','0','1','1','0','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
