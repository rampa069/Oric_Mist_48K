
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"fd",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"f4",x"fd",x"c2"),
    18 => (x"48",x"cc",x"e5",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"c9",x"e5",x"c2",x"87"),
    25 => (x"c5",x"e5",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e9",x"c1",x"87",x"f7"),
    29 => (x"e5",x"c2",x"87",x"f1"),
    30 => (x"e5",x"c2",x"4d",x"c9"),
    31 => (x"ad",x"74",x"4c",x"c9"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"cf",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"df",x"4c",x"87",x"c9"),
    69 => (x"88",x"74",x"9c",x"98"),
    70 => (x"26",x"87",x"ec",x"02"),
    71 => (x"26",x"4b",x"26",x"4a"),
    72 => (x"1e",x"4f",x"26",x"4c"),
    73 => (x"73",x"81",x"48",x"73"),
    74 => (x"87",x"c5",x"02",x"a9"),
    75 => (x"f6",x"05",x"53",x"12"),
    76 => (x"1e",x"4f",x"26",x"87"),
    77 => (x"4a",x"71",x"1e",x"73"),
    78 => (x"49",x"4b",x"66",x"c8"),
    79 => (x"99",x"71",x"8b",x"c1"),
    80 => (x"12",x"87",x"cf",x"02"),
    81 => (x"08",x"d4",x"ff",x"48"),
    82 => (x"c1",x"49",x"73",x"78"),
    83 => (x"05",x"99",x"71",x"8b"),
    84 => (x"4b",x"26",x"87",x"f1"),
    85 => (x"5e",x"0e",x"4f",x"26"),
    86 => (x"71",x"0e",x"5c",x"5b"),
    87 => (x"4c",x"d4",x"ff",x"4a"),
    88 => (x"49",x"4b",x"66",x"cc"),
    89 => (x"99",x"71",x"8b",x"c1"),
    90 => (x"c3",x"87",x"ce",x"02"),
    91 => (x"52",x"6c",x"7c",x"ff"),
    92 => (x"8b",x"c1",x"49",x"73"),
    93 => (x"f2",x"05",x"99",x"71"),
    94 => (x"26",x"4c",x"26",x"87"),
    95 => (x"1e",x"4f",x"26",x"4b"),
    96 => (x"d4",x"ff",x"1e",x"73"),
    97 => (x"7b",x"ff",x"c3",x"4b"),
    98 => (x"ff",x"c3",x"4a",x"6b"),
    99 => (x"c8",x"49",x"6b",x"7b"),
   100 => (x"c3",x"b1",x"72",x"32"),
   101 => (x"4a",x"6b",x"7b",x"ff"),
   102 => (x"b2",x"71",x"31",x"c8"),
   103 => (x"6b",x"7b",x"ff",x"c3"),
   104 => (x"72",x"32",x"c8",x"49"),
   105 => (x"26",x"48",x"71",x"b1"),
   106 => (x"0e",x"4f",x"26",x"4b"),
   107 => (x"5d",x"5c",x"5b",x"5e"),
   108 => (x"ff",x"4d",x"71",x"0e"),
   109 => (x"48",x"75",x"4c",x"d4"),
   110 => (x"70",x"98",x"ff",x"c3"),
   111 => (x"cc",x"e5",x"c2",x"7c"),
   112 => (x"87",x"c8",x"05",x"bf"),
   113 => (x"c9",x"48",x"66",x"d0"),
   114 => (x"58",x"a6",x"d4",x"30"),
   115 => (x"d8",x"49",x"66",x"d0"),
   116 => (x"c3",x"48",x"71",x"29"),
   117 => (x"7c",x"70",x"98",x"ff"),
   118 => (x"d0",x"49",x"66",x"d0"),
   119 => (x"c3",x"48",x"71",x"29"),
   120 => (x"7c",x"70",x"98",x"ff"),
   121 => (x"c8",x"49",x"66",x"d0"),
   122 => (x"c3",x"48",x"71",x"29"),
   123 => (x"7c",x"70",x"98",x"ff"),
   124 => (x"c3",x"48",x"66",x"d0"),
   125 => (x"7c",x"70",x"98",x"ff"),
   126 => (x"29",x"d0",x"49",x"75"),
   127 => (x"ff",x"c3",x"48",x"71"),
   128 => (x"6c",x"7c",x"70",x"98"),
   129 => (x"ff",x"f0",x"c9",x"4b"),
   130 => (x"ab",x"ff",x"c3",x"4a"),
   131 => (x"49",x"87",x"cf",x"05"),
   132 => (x"4b",x"6c",x"7c",x"71"),
   133 => (x"c5",x"02",x"8a",x"c1"),
   134 => (x"02",x"ab",x"71",x"87"),
   135 => (x"48",x"73",x"87",x"f2"),
   136 => (x"4c",x"26",x"4d",x"26"),
   137 => (x"4f",x"26",x"4b",x"26"),
   138 => (x"ff",x"49",x"c0",x"1e"),
   139 => (x"ff",x"c3",x"48",x"d4"),
   140 => (x"c3",x"81",x"c1",x"78"),
   141 => (x"04",x"a9",x"b7",x"c8"),
   142 => (x"4f",x"26",x"87",x"f1"),
   143 => (x"5c",x"5b",x"5e",x"0e"),
   144 => (x"ff",x"c0",x"0e",x"5d"),
   145 => (x"4d",x"f7",x"c1",x"f0"),
   146 => (x"c0",x"c0",x"c0",x"c1"),
   147 => (x"ff",x"4b",x"c0",x"c0"),
   148 => (x"f8",x"c4",x"87",x"d6"),
   149 => (x"1e",x"c0",x"4c",x"df"),
   150 => (x"ce",x"fd",x"49",x"75"),
   151 => (x"c1",x"86",x"c4",x"87"),
   152 => (x"e5",x"c0",x"05",x"a8"),
   153 => (x"48",x"d4",x"ff",x"87"),
   154 => (x"73",x"78",x"ff",x"c3"),
   155 => (x"f0",x"e1",x"c0",x"1e"),
   156 => (x"fc",x"49",x"e9",x"c1"),
   157 => (x"86",x"c4",x"87",x"f5"),
   158 => (x"ca",x"05",x"98",x"70"),
   159 => (x"48",x"d4",x"ff",x"87"),
   160 => (x"c1",x"78",x"ff",x"c3"),
   161 => (x"fe",x"87",x"cb",x"48"),
   162 => (x"8c",x"c1",x"87",x"de"),
   163 => (x"87",x"c6",x"ff",x"05"),
   164 => (x"4d",x"26",x"48",x"c0"),
   165 => (x"4b",x"26",x"4c",x"26"),
   166 => (x"5e",x"0e",x"4f",x"26"),
   167 => (x"c0",x"0e",x"5c",x"5b"),
   168 => (x"c1",x"c1",x"f0",x"ff"),
   169 => (x"48",x"d4",x"ff",x"4c"),
   170 => (x"cb",x"78",x"ff",x"c3"),
   171 => (x"f6",x"f7",x"49",x"dc"),
   172 => (x"c0",x"4b",x"d3",x"87"),
   173 => (x"fb",x"49",x"74",x"1e"),
   174 => (x"86",x"c4",x"87",x"f1"),
   175 => (x"ca",x"05",x"98",x"70"),
   176 => (x"48",x"d4",x"ff",x"87"),
   177 => (x"c1",x"78",x"ff",x"c3"),
   178 => (x"fd",x"87",x"cb",x"48"),
   179 => (x"8b",x"c1",x"87",x"da"),
   180 => (x"87",x"df",x"ff",x"05"),
   181 => (x"4c",x"26",x"48",x"c0"),
   182 => (x"4f",x"26",x"4b",x"26"),
   183 => (x"00",x"44",x"4d",x"43"),
   184 => (x"43",x"48",x"44",x"53"),
   185 => (x"69",x"61",x"66",x"20"),
   186 => (x"00",x"0a",x"21",x"6c"),
   187 => (x"52",x"52",x"45",x"49"),
   188 => (x"00",x"00",x"00",x"00"),
   189 => (x"00",x"49",x"50",x"53"),
   190 => (x"74",x"69",x"72",x"57"),
   191 => (x"61",x"66",x"20",x"65"),
   192 => (x"64",x"65",x"6c",x"69"),
   193 => (x"5e",x"0e",x"00",x"0a"),
   194 => (x"0e",x"5d",x"5c",x"5b"),
   195 => (x"ff",x"4d",x"ff",x"c3"),
   196 => (x"d3",x"fc",x"4b",x"d4"),
   197 => (x"1e",x"ea",x"c6",x"87"),
   198 => (x"c1",x"f0",x"e1",x"c0"),
   199 => (x"ca",x"fa",x"49",x"c8"),
   200 => (x"c1",x"86",x"c4",x"87"),
   201 => (x"87",x"c8",x"02",x"a8"),
   202 => (x"c0",x"87",x"ef",x"fd"),
   203 => (x"87",x"e8",x"c1",x"48"),
   204 => (x"70",x"87",x"cc",x"f9"),
   205 => (x"ff",x"ff",x"cf",x"49"),
   206 => (x"a9",x"ea",x"c6",x"99"),
   207 => (x"fd",x"87",x"c8",x"02"),
   208 => (x"48",x"c0",x"87",x"d8"),
   209 => (x"75",x"87",x"d1",x"c1"),
   210 => (x"4c",x"f1",x"c0",x"7b"),
   211 => (x"70",x"87",x"ed",x"fb"),
   212 => (x"ec",x"c0",x"02",x"98"),
   213 => (x"c0",x"1e",x"c0",x"87"),
   214 => (x"fa",x"c1",x"f0",x"ff"),
   215 => (x"87",x"cb",x"f9",x"49"),
   216 => (x"98",x"70",x"86",x"c4"),
   217 => (x"75",x"87",x"da",x"05"),
   218 => (x"75",x"49",x"6b",x"7b"),
   219 => (x"75",x"7b",x"75",x"7b"),
   220 => (x"c1",x"7b",x"75",x"7b"),
   221 => (x"c4",x"02",x"99",x"c0"),
   222 => (x"db",x"48",x"c1",x"87"),
   223 => (x"d7",x"48",x"c0",x"87"),
   224 => (x"05",x"ac",x"c2",x"87"),
   225 => (x"e0",x"cb",x"87",x"ca"),
   226 => (x"87",x"db",x"f4",x"49"),
   227 => (x"87",x"c8",x"48",x"c0"),
   228 => (x"fe",x"05",x"8c",x"c1"),
   229 => (x"48",x"c0",x"87",x"f6"),
   230 => (x"4c",x"26",x"4d",x"26"),
   231 => (x"4f",x"26",x"4b",x"26"),
   232 => (x"5c",x"5b",x"5e",x"0e"),
   233 => (x"d0",x"ff",x"0e",x"5d"),
   234 => (x"d0",x"e5",x"c0",x"4d"),
   235 => (x"c2",x"4c",x"c0",x"c1"),
   236 => (x"c1",x"48",x"cc",x"e5"),
   237 => (x"49",x"f4",x"cb",x"78"),
   238 => (x"c7",x"87",x"ec",x"f3"),
   239 => (x"f9",x"7d",x"c2",x"4b"),
   240 => (x"7d",x"c3",x"87",x"e6"),
   241 => (x"49",x"74",x"1e",x"c0"),
   242 => (x"c4",x"87",x"e0",x"f7"),
   243 => (x"05",x"a8",x"c1",x"86"),
   244 => (x"c2",x"4b",x"87",x"c1"),
   245 => (x"87",x"cb",x"05",x"ab"),
   246 => (x"f3",x"49",x"ec",x"cb"),
   247 => (x"48",x"c0",x"87",x"c9"),
   248 => (x"c1",x"87",x"f6",x"c0"),
   249 => (x"d4",x"ff",x"05",x"8b"),
   250 => (x"87",x"da",x"fc",x"87"),
   251 => (x"58",x"d0",x"e5",x"c2"),
   252 => (x"cd",x"05",x"98",x"70"),
   253 => (x"c0",x"1e",x"c1",x"87"),
   254 => (x"d0",x"c1",x"f0",x"ff"),
   255 => (x"87",x"eb",x"f6",x"49"),
   256 => (x"d4",x"ff",x"86",x"c4"),
   257 => (x"78",x"ff",x"c3",x"48"),
   258 => (x"c2",x"87",x"ee",x"c4"),
   259 => (x"c2",x"58",x"d4",x"e5"),
   260 => (x"48",x"d4",x"ff",x"7d"),
   261 => (x"c1",x"78",x"ff",x"c3"),
   262 => (x"26",x"4d",x"26",x"48"),
   263 => (x"26",x"4b",x"26",x"4c"),
   264 => (x"5b",x"5e",x"0e",x"4f"),
   265 => (x"71",x"0e",x"5d",x"5c"),
   266 => (x"4c",x"ff",x"c3",x"4d"),
   267 => (x"74",x"4b",x"d4",x"ff"),
   268 => (x"48",x"d0",x"ff",x"7b"),
   269 => (x"74",x"78",x"c3",x"c4"),
   270 => (x"c0",x"1e",x"75",x"7b"),
   271 => (x"d8",x"c1",x"f0",x"ff"),
   272 => (x"87",x"e7",x"f5",x"49"),
   273 => (x"98",x"70",x"86",x"c4"),
   274 => (x"cb",x"87",x"cb",x"02"),
   275 => (x"d6",x"f1",x"49",x"f8"),
   276 => (x"c0",x"48",x"c1",x"87"),
   277 => (x"7b",x"74",x"87",x"ee"),
   278 => (x"c8",x"7b",x"fe",x"c3"),
   279 => (x"66",x"d4",x"1e",x"c0"),
   280 => (x"87",x"cf",x"f3",x"49"),
   281 => (x"7b",x"74",x"86",x"c4"),
   282 => (x"7b",x"74",x"7b",x"74"),
   283 => (x"4a",x"e0",x"da",x"d8"),
   284 => (x"05",x"6b",x"7b",x"74"),
   285 => (x"8a",x"c1",x"87",x"c5"),
   286 => (x"74",x"87",x"f5",x"05"),
   287 => (x"48",x"d0",x"ff",x"7b"),
   288 => (x"48",x"c0",x"78",x"c2"),
   289 => (x"4c",x"26",x"4d",x"26"),
   290 => (x"4f",x"26",x"4b",x"26"),
   291 => (x"5c",x"5b",x"5e",x"0e"),
   292 => (x"86",x"fc",x"0e",x"5d"),
   293 => (x"d4",x"ff",x"4b",x"71"),
   294 => (x"c5",x"7e",x"c0",x"4c"),
   295 => (x"4a",x"df",x"cd",x"ee"),
   296 => (x"6c",x"7c",x"ff",x"c3"),
   297 => (x"a8",x"fe",x"c3",x"48"),
   298 => (x"87",x"f8",x"c0",x"05"),
   299 => (x"9b",x"73",x"4d",x"74"),
   300 => (x"d4",x"87",x"cc",x"02"),
   301 => (x"49",x"73",x"1e",x"66"),
   302 => (x"c4",x"87",x"db",x"f2"),
   303 => (x"ff",x"87",x"d4",x"86"),
   304 => (x"d1",x"c4",x"48",x"d0"),
   305 => (x"4a",x"66",x"d4",x"78"),
   306 => (x"c1",x"7d",x"ff",x"c3"),
   307 => (x"87",x"f8",x"05",x"8a"),
   308 => (x"c3",x"5a",x"a6",x"d8"),
   309 => (x"73",x"7c",x"7c",x"ff"),
   310 => (x"87",x"c5",x"05",x"9b"),
   311 => (x"d0",x"48",x"d0",x"ff"),
   312 => (x"7e",x"4a",x"c1",x"78"),
   313 => (x"fe",x"05",x"8a",x"c1"),
   314 => (x"48",x"6e",x"87",x"f6"),
   315 => (x"4d",x"26",x"8e",x"fc"),
   316 => (x"4b",x"26",x"4c",x"26"),
   317 => (x"73",x"1e",x"4f",x"26"),
   318 => (x"c0",x"4a",x"71",x"1e"),
   319 => (x"48",x"d4",x"ff",x"4b"),
   320 => (x"ff",x"78",x"ff",x"c3"),
   321 => (x"c3",x"c4",x"48",x"d0"),
   322 => (x"48",x"d4",x"ff",x"78"),
   323 => (x"72",x"78",x"ff",x"c3"),
   324 => (x"f0",x"ff",x"c0",x"1e"),
   325 => (x"f2",x"49",x"d1",x"c1"),
   326 => (x"86",x"c4",x"87",x"d1"),
   327 => (x"d2",x"05",x"98",x"70"),
   328 => (x"1e",x"c0",x"c8",x"87"),
   329 => (x"fd",x"49",x"66",x"cc"),
   330 => (x"86",x"c4",x"87",x"e2"),
   331 => (x"d0",x"ff",x"4b",x"70"),
   332 => (x"73",x"78",x"c2",x"48"),
   333 => (x"26",x"4b",x"26",x"48"),
   334 => (x"5b",x"5e",x"0e",x"4f"),
   335 => (x"c0",x"0e",x"5d",x"5c"),
   336 => (x"f0",x"ff",x"c0",x"1e"),
   337 => (x"f1",x"49",x"c9",x"c1"),
   338 => (x"1e",x"d2",x"87",x"e1"),
   339 => (x"49",x"dc",x"e5",x"c2"),
   340 => (x"c8",x"87",x"f9",x"fc"),
   341 => (x"c1",x"4c",x"c0",x"86"),
   342 => (x"ac",x"b7",x"d2",x"84"),
   343 => (x"c2",x"87",x"f8",x"04"),
   344 => (x"bf",x"97",x"dc",x"e5"),
   345 => (x"99",x"c0",x"c3",x"49"),
   346 => (x"05",x"a9",x"c0",x"c1"),
   347 => (x"c2",x"87",x"e7",x"c0"),
   348 => (x"bf",x"97",x"e3",x"e5"),
   349 => (x"c2",x"31",x"d0",x"49"),
   350 => (x"bf",x"97",x"e4",x"e5"),
   351 => (x"72",x"32",x"c8",x"4a"),
   352 => (x"e5",x"e5",x"c2",x"b1"),
   353 => (x"b1",x"4a",x"bf",x"97"),
   354 => (x"ff",x"cf",x"4c",x"71"),
   355 => (x"c1",x"9c",x"ff",x"ff"),
   356 => (x"c1",x"34",x"ca",x"84"),
   357 => (x"e5",x"c2",x"87",x"e7"),
   358 => (x"49",x"bf",x"97",x"e5"),
   359 => (x"99",x"c6",x"31",x"c1"),
   360 => (x"97",x"e6",x"e5",x"c2"),
   361 => (x"b7",x"c7",x"4a",x"bf"),
   362 => (x"c2",x"b1",x"72",x"2a"),
   363 => (x"bf",x"97",x"e1",x"e5"),
   364 => (x"9d",x"cf",x"4d",x"4a"),
   365 => (x"97",x"e2",x"e5",x"c2"),
   366 => (x"9a",x"c3",x"4a",x"bf"),
   367 => (x"e5",x"c2",x"32",x"ca"),
   368 => (x"4b",x"bf",x"97",x"e3"),
   369 => (x"b2",x"73",x"33",x"c2"),
   370 => (x"97",x"e4",x"e5",x"c2"),
   371 => (x"c0",x"c3",x"4b",x"bf"),
   372 => (x"2b",x"b7",x"c6",x"9b"),
   373 => (x"81",x"c2",x"b2",x"73"),
   374 => (x"30",x"71",x"48",x"c1"),
   375 => (x"48",x"c1",x"49",x"70"),
   376 => (x"4d",x"70",x"30",x"75"),
   377 => (x"84",x"c1",x"4c",x"72"),
   378 => (x"c0",x"c8",x"94",x"71"),
   379 => (x"cc",x"06",x"ad",x"b7"),
   380 => (x"b7",x"34",x"c1",x"87"),
   381 => (x"b7",x"c0",x"c8",x"2d"),
   382 => (x"f4",x"ff",x"01",x"ad"),
   383 => (x"26",x"48",x"74",x"87"),
   384 => (x"26",x"4c",x"26",x"4d"),
   385 => (x"0e",x"4f",x"26",x"4b"),
   386 => (x"5d",x"5c",x"5b",x"5e"),
   387 => (x"c2",x"86",x"fc",x"0e"),
   388 => (x"c0",x"48",x"c4",x"ee"),
   389 => (x"fc",x"e5",x"c2",x"78"),
   390 => (x"fb",x"49",x"c0",x"1e"),
   391 => (x"86",x"c4",x"87",x"d8"),
   392 => (x"c5",x"05",x"98",x"70"),
   393 => (x"c9",x"48",x"c0",x"87"),
   394 => (x"4d",x"c0",x"87",x"d2"),
   395 => (x"48",x"c0",x"f3",x"c2"),
   396 => (x"e6",x"c2",x"78",x"c1"),
   397 => (x"e2",x"c0",x"4a",x"f2"),
   398 => (x"4b",x"c8",x"49",x"d4"),
   399 => (x"70",x"87",x"e7",x"ea"),
   400 => (x"87",x"c6",x"05",x"98"),
   401 => (x"48",x"c0",x"f3",x"c2"),
   402 => (x"e7",x"c2",x"78",x"c0"),
   403 => (x"e2",x"c0",x"4a",x"ce"),
   404 => (x"4b",x"c8",x"49",x"e0"),
   405 => (x"70",x"87",x"cf",x"ea"),
   406 => (x"87",x"c6",x"05",x"98"),
   407 => (x"48",x"c0",x"f3",x"c2"),
   408 => (x"f3",x"c2",x"78",x"c0"),
   409 => (x"c0",x"02",x"bf",x"c0"),
   410 => (x"ed",x"c2",x"87",x"fd"),
   411 => (x"c2",x"4d",x"bf",x"c2"),
   412 => (x"bf",x"9f",x"fa",x"ed"),
   413 => (x"d6",x"c5",x"48",x"7e"),
   414 => (x"c7",x"05",x"a8",x"ea"),
   415 => (x"c2",x"ed",x"c2",x"87"),
   416 => (x"87",x"ce",x"4d",x"bf"),
   417 => (x"e9",x"ca",x"48",x"6e"),
   418 => (x"c5",x"02",x"a8",x"d5"),
   419 => (x"c7",x"48",x"c0",x"87"),
   420 => (x"e5",x"c2",x"87",x"ea"),
   421 => (x"49",x"75",x"1e",x"fc"),
   422 => (x"c4",x"87",x"db",x"f9"),
   423 => (x"05",x"98",x"70",x"86"),
   424 => (x"48",x"c0",x"87",x"c5"),
   425 => (x"c2",x"87",x"d5",x"c7"),
   426 => (x"c0",x"4a",x"ce",x"e7"),
   427 => (x"c8",x"49",x"ec",x"e2"),
   428 => (x"87",x"f2",x"e8",x"4b"),
   429 => (x"c8",x"05",x"98",x"70"),
   430 => (x"c4",x"ee",x"c2",x"87"),
   431 => (x"d8",x"78",x"c1",x"48"),
   432 => (x"f2",x"e6",x"c2",x"87"),
   433 => (x"f8",x"e2",x"c0",x"4a"),
   434 => (x"e8",x"4b",x"c8",x"49"),
   435 => (x"98",x"70",x"87",x"d8"),
   436 => (x"87",x"c5",x"c0",x"02"),
   437 => (x"e3",x"c6",x"48",x"c0"),
   438 => (x"fa",x"ed",x"c2",x"87"),
   439 => (x"c1",x"49",x"bf",x"97"),
   440 => (x"c0",x"05",x"a9",x"d5"),
   441 => (x"ed",x"c2",x"87",x"cd"),
   442 => (x"49",x"bf",x"97",x"fb"),
   443 => (x"02",x"a9",x"ea",x"c2"),
   444 => (x"c0",x"87",x"c5",x"c0"),
   445 => (x"87",x"c4",x"c6",x"48"),
   446 => (x"97",x"fc",x"e5",x"c2"),
   447 => (x"c3",x"48",x"7e",x"bf"),
   448 => (x"c0",x"02",x"a8",x"e9"),
   449 => (x"48",x"6e",x"87",x"ce"),
   450 => (x"02",x"a8",x"eb",x"c3"),
   451 => (x"c0",x"87",x"c5",x"c0"),
   452 => (x"87",x"e8",x"c5",x"48"),
   453 => (x"97",x"c7",x"e6",x"c2"),
   454 => (x"05",x"99",x"49",x"bf"),
   455 => (x"c2",x"87",x"cc",x"c0"),
   456 => (x"bf",x"97",x"c8",x"e6"),
   457 => (x"02",x"a9",x"c2",x"49"),
   458 => (x"c0",x"87",x"c5",x"c0"),
   459 => (x"87",x"cc",x"c5",x"48"),
   460 => (x"97",x"c9",x"e6",x"c2"),
   461 => (x"ee",x"c2",x"48",x"bf"),
   462 => (x"4c",x"70",x"58",x"c0"),
   463 => (x"c2",x"88",x"c1",x"48"),
   464 => (x"c2",x"58",x"c4",x"ee"),
   465 => (x"bf",x"97",x"ca",x"e6"),
   466 => (x"c2",x"81",x"75",x"49"),
   467 => (x"bf",x"97",x"cb",x"e6"),
   468 => (x"72",x"32",x"c8",x"4a"),
   469 => (x"f2",x"c2",x"7e",x"a1"),
   470 => (x"78",x"6e",x"48",x"dc"),
   471 => (x"97",x"cc",x"e6",x"c2"),
   472 => (x"f2",x"c2",x"48",x"bf"),
   473 => (x"ee",x"c2",x"58",x"f4"),
   474 => (x"c2",x"02",x"bf",x"c4"),
   475 => (x"e7",x"c2",x"87",x"d3"),
   476 => (x"e2",x"c0",x"4a",x"ce"),
   477 => (x"4b",x"c8",x"49",x"c8"),
   478 => (x"70",x"87",x"eb",x"e5"),
   479 => (x"c5",x"c0",x"02",x"98"),
   480 => (x"c3",x"48",x"c0",x"87"),
   481 => (x"ed",x"c2",x"87",x"f6"),
   482 => (x"c2",x"4c",x"bf",x"fc"),
   483 => (x"c2",x"5c",x"f0",x"f2"),
   484 => (x"bf",x"97",x"e1",x"e6"),
   485 => (x"c2",x"31",x"c8",x"49"),
   486 => (x"bf",x"97",x"e0",x"e6"),
   487 => (x"c2",x"49",x"a1",x"4a"),
   488 => (x"bf",x"97",x"e2",x"e6"),
   489 => (x"72",x"32",x"d0",x"4a"),
   490 => (x"e6",x"c2",x"49",x"a1"),
   491 => (x"4a",x"bf",x"97",x"e3"),
   492 => (x"a1",x"72",x"32",x"d8"),
   493 => (x"f8",x"f2",x"c2",x"49"),
   494 => (x"f0",x"f2",x"c2",x"59"),
   495 => (x"f2",x"c2",x"91",x"bf"),
   496 => (x"c2",x"81",x"bf",x"dc"),
   497 => (x"c2",x"59",x"e4",x"f2"),
   498 => (x"bf",x"97",x"e9",x"e6"),
   499 => (x"c2",x"32",x"c8",x"4a"),
   500 => (x"bf",x"97",x"e8",x"e6"),
   501 => (x"c2",x"4a",x"a2",x"4b"),
   502 => (x"bf",x"97",x"ea",x"e6"),
   503 => (x"73",x"33",x"d0",x"4b"),
   504 => (x"e6",x"c2",x"4a",x"a2"),
   505 => (x"4b",x"bf",x"97",x"eb"),
   506 => (x"33",x"d8",x"9b",x"cf"),
   507 => (x"c2",x"4a",x"a2",x"73"),
   508 => (x"c2",x"5a",x"e8",x"f2"),
   509 => (x"c2",x"92",x"74",x"8a"),
   510 => (x"72",x"48",x"e8",x"f2"),
   511 => (x"c7",x"c1",x"78",x"a1"),
   512 => (x"ce",x"e6",x"c2",x"87"),
   513 => (x"c8",x"49",x"bf",x"97"),
   514 => (x"cd",x"e6",x"c2",x"31"),
   515 => (x"a1",x"4a",x"bf",x"97"),
   516 => (x"c7",x"31",x"c5",x"49"),
   517 => (x"29",x"c9",x"81",x"ff"),
   518 => (x"59",x"f0",x"f2",x"c2"),
   519 => (x"97",x"d3",x"e6",x"c2"),
   520 => (x"32",x"c8",x"4a",x"bf"),
   521 => (x"97",x"d2",x"e6",x"c2"),
   522 => (x"4a",x"a2",x"4b",x"bf"),
   523 => (x"5a",x"f8",x"f2",x"c2"),
   524 => (x"bf",x"f0",x"f2",x"c2"),
   525 => (x"c2",x"82",x"6e",x"92"),
   526 => (x"c2",x"5a",x"ec",x"f2"),
   527 => (x"c0",x"48",x"e4",x"f2"),
   528 => (x"e0",x"f2",x"c2",x"78"),
   529 => (x"78",x"a1",x"72",x"48"),
   530 => (x"48",x"f8",x"f2",x"c2"),
   531 => (x"bf",x"e4",x"f2",x"c2"),
   532 => (x"fc",x"f2",x"c2",x"78"),
   533 => (x"e8",x"f2",x"c2",x"48"),
   534 => (x"ee",x"c2",x"78",x"bf"),
   535 => (x"c0",x"02",x"bf",x"c4"),
   536 => (x"48",x"74",x"87",x"c9"),
   537 => (x"7e",x"70",x"30",x"c4"),
   538 => (x"c2",x"87",x"c9",x"c0"),
   539 => (x"48",x"bf",x"ec",x"f2"),
   540 => (x"7e",x"70",x"30",x"c4"),
   541 => (x"48",x"c8",x"ee",x"c2"),
   542 => (x"48",x"c1",x"78",x"6e"),
   543 => (x"4d",x"26",x"8e",x"fc"),
   544 => (x"4b",x"26",x"4c",x"26"),
   545 => (x"00",x"00",x"4f",x"26"),
   546 => (x"33",x"54",x"41",x"46"),
   547 => (x"20",x"20",x"20",x"32"),
   548 => (x"00",x"00",x"00",x"00"),
   549 => (x"31",x"54",x"41",x"46"),
   550 => (x"20",x"20",x"20",x"36"),
   551 => (x"00",x"00",x"00",x"00"),
   552 => (x"33",x"54",x"41",x"46"),
   553 => (x"20",x"20",x"20",x"32"),
   554 => (x"00",x"00",x"00",x"00"),
   555 => (x"33",x"54",x"41",x"46"),
   556 => (x"20",x"20",x"20",x"32"),
   557 => (x"00",x"00",x"00",x"00"),
   558 => (x"31",x"54",x"41",x"46"),
   559 => (x"20",x"20",x"20",x"36"),
   560 => (x"5b",x"5e",x"0e",x"00"),
   561 => (x"71",x"0e",x"5d",x"5c"),
   562 => (x"c4",x"ee",x"c2",x"4a"),
   563 => (x"87",x"cb",x"02",x"bf"),
   564 => (x"2b",x"c7",x"4b",x"72"),
   565 => (x"ff",x"c1",x"4d",x"72"),
   566 => (x"72",x"87",x"c9",x"9d"),
   567 => (x"72",x"2b",x"c8",x"4b"),
   568 => (x"9d",x"ff",x"c3",x"4d"),
   569 => (x"bf",x"dc",x"f2",x"c2"),
   570 => (x"cc",x"fa",x"c0",x"83"),
   571 => (x"d9",x"02",x"ab",x"bf"),
   572 => (x"d0",x"fa",x"c0",x"87"),
   573 => (x"fc",x"e5",x"c2",x"5b"),
   574 => (x"ef",x"49",x"73",x"1e"),
   575 => (x"86",x"c4",x"87",x"f8"),
   576 => (x"c5",x"05",x"98",x"70"),
   577 => (x"c0",x"48",x"c0",x"87"),
   578 => (x"ee",x"c2",x"87",x"e6"),
   579 => (x"d2",x"02",x"bf",x"c4"),
   580 => (x"c4",x"49",x"75",x"87"),
   581 => (x"fc",x"e5",x"c2",x"91"),
   582 => (x"cf",x"4c",x"69",x"81"),
   583 => (x"ff",x"ff",x"ff",x"ff"),
   584 => (x"75",x"87",x"cb",x"9c"),
   585 => (x"c2",x"91",x"c2",x"49"),
   586 => (x"9f",x"81",x"fc",x"e5"),
   587 => (x"48",x"74",x"4c",x"69"),
   588 => (x"4c",x"26",x"4d",x"26"),
   589 => (x"4f",x"26",x"4b",x"26"),
   590 => (x"5c",x"5b",x"5e",x"0e"),
   591 => (x"86",x"f4",x"0e",x"5d"),
   592 => (x"c4",x"59",x"a6",x"c8"),
   593 => (x"80",x"c8",x"48",x"66"),
   594 => (x"c0",x"48",x"7e",x"70"),
   595 => (x"49",x"c1",x"1e",x"78"),
   596 => (x"87",x"fd",x"cc",x"49"),
   597 => (x"4c",x"70",x"86",x"c4"),
   598 => (x"fc",x"c0",x"02",x"9c"),
   599 => (x"cc",x"ee",x"c2",x"87"),
   600 => (x"49",x"66",x"dc",x"4a"),
   601 => (x"87",x"e3",x"dd",x"ff"),
   602 => (x"c0",x"02",x"98",x"70"),
   603 => (x"4a",x"74",x"87",x"eb"),
   604 => (x"cb",x"49",x"66",x"dc"),
   605 => (x"c7",x"de",x"ff",x"4b"),
   606 => (x"02",x"98",x"70",x"87"),
   607 => (x"1e",x"c0",x"87",x"db"),
   608 => (x"c4",x"02",x"9c",x"74"),
   609 => (x"c2",x"4d",x"c0",x"87"),
   610 => (x"75",x"4d",x"c1",x"87"),
   611 => (x"87",x"c1",x"cc",x"49"),
   612 => (x"4c",x"70",x"86",x"c4"),
   613 => (x"c4",x"ff",x"05",x"9c"),
   614 => (x"02",x"9c",x"74",x"87"),
   615 => (x"dc",x"87",x"f4",x"c1"),
   616 => (x"48",x"6e",x"49",x"a4"),
   617 => (x"a4",x"da",x"78",x"69"),
   618 => (x"4d",x"66",x"c4",x"49"),
   619 => (x"69",x"9f",x"85",x"c4"),
   620 => (x"c4",x"ee",x"c2",x"7d"),
   621 => (x"87",x"d2",x"02",x"bf"),
   622 => (x"9f",x"49",x"a4",x"d4"),
   623 => (x"ff",x"c0",x"49",x"69"),
   624 => (x"48",x"71",x"99",x"ff"),
   625 => (x"7e",x"70",x"30",x"d0"),
   626 => (x"7e",x"c0",x"87",x"c2"),
   627 => (x"6d",x"48",x"49",x"6e"),
   628 => (x"c4",x"7d",x"70",x"80"),
   629 => (x"78",x"c0",x"48",x"66"),
   630 => (x"cc",x"49",x"66",x"c4"),
   631 => (x"c4",x"79",x"6d",x"81"),
   632 => (x"81",x"d0",x"49",x"66"),
   633 => (x"a6",x"c8",x"79",x"c0"),
   634 => (x"c8",x"78",x"c0",x"48"),
   635 => (x"66",x"c4",x"4c",x"66"),
   636 => (x"74",x"82",x"d4",x"4a"),
   637 => (x"72",x"91",x"c8",x"49"),
   638 => (x"41",x"c0",x"49",x"a1"),
   639 => (x"84",x"c1",x"79",x"6d"),
   640 => (x"04",x"ac",x"b7",x"c6"),
   641 => (x"c4",x"87",x"e7",x"ff"),
   642 => (x"c4",x"c1",x"49",x"66"),
   643 => (x"c1",x"79",x"c0",x"81"),
   644 => (x"c0",x"87",x"c2",x"48"),
   645 => (x"26",x"8e",x"f4",x"48"),
   646 => (x"26",x"4c",x"26",x"4d"),
   647 => (x"0e",x"4f",x"26",x"4b"),
   648 => (x"5d",x"5c",x"5b",x"5e"),
   649 => (x"d0",x"4c",x"71",x"0e"),
   650 => (x"49",x"6c",x"4d",x"66"),
   651 => (x"c2",x"b9",x"75",x"85"),
   652 => (x"4a",x"bf",x"c0",x"ee"),
   653 => (x"99",x"72",x"ba",x"ff"),
   654 => (x"c0",x"02",x"99",x"71"),
   655 => (x"a4",x"c4",x"87",x"e4"),
   656 => (x"f9",x"49",x"6b",x"4b"),
   657 => (x"7b",x"70",x"87",x"fb"),
   658 => (x"bf",x"fc",x"ed",x"c2"),
   659 => (x"71",x"81",x"6c",x"49"),
   660 => (x"c2",x"b9",x"75",x"7c"),
   661 => (x"4a",x"bf",x"c0",x"ee"),
   662 => (x"99",x"72",x"ba",x"ff"),
   663 => (x"ff",x"05",x"99",x"71"),
   664 => (x"7c",x"75",x"87",x"dc"),
   665 => (x"4c",x"26",x"4d",x"26"),
   666 => (x"4f",x"26",x"4b",x"26"),
   667 => (x"71",x"1e",x"73",x"1e"),
   668 => (x"e0",x"f2",x"c2",x"4b"),
   669 => (x"a3",x"c4",x"49",x"bf"),
   670 => (x"c2",x"4a",x"6a",x"4a"),
   671 => (x"fc",x"ed",x"c2",x"8a"),
   672 => (x"a1",x"72",x"92",x"bf"),
   673 => (x"c0",x"ee",x"c2",x"49"),
   674 => (x"9a",x"6b",x"4a",x"bf"),
   675 => (x"c0",x"49",x"a1",x"72"),
   676 => (x"c8",x"59",x"d0",x"fa"),
   677 => (x"e9",x"71",x"1e",x"66"),
   678 => (x"86",x"c4",x"87",x"dc"),
   679 => (x"c4",x"05",x"98",x"70"),
   680 => (x"c2",x"48",x"c0",x"87"),
   681 => (x"26",x"48",x"c1",x"87"),
   682 => (x"1e",x"4f",x"26",x"4b"),
   683 => (x"4b",x"71",x"1e",x"73"),
   684 => (x"bf",x"e0",x"f2",x"c2"),
   685 => (x"4a",x"a3",x"c4",x"49"),
   686 => (x"8a",x"c2",x"4a",x"6a"),
   687 => (x"bf",x"fc",x"ed",x"c2"),
   688 => (x"49",x"a1",x"72",x"92"),
   689 => (x"bf",x"c0",x"ee",x"c2"),
   690 => (x"72",x"9a",x"6b",x"4a"),
   691 => (x"fa",x"c0",x"49",x"a1"),
   692 => (x"66",x"c8",x"59",x"d0"),
   693 => (x"c8",x"e5",x"71",x"1e"),
   694 => (x"70",x"86",x"c4",x"87"),
   695 => (x"87",x"c4",x"05",x"98"),
   696 => (x"87",x"c2",x"48",x"c0"),
   697 => (x"4b",x"26",x"48",x"c1"),
   698 => (x"5e",x"0e",x"4f",x"26"),
   699 => (x"0e",x"5d",x"5c",x"5b"),
   700 => (x"4b",x"71",x"86",x"e4"),
   701 => (x"48",x"66",x"ec",x"c0"),
   702 => (x"a6",x"cc",x"28",x"c9"),
   703 => (x"c0",x"ee",x"c2",x"58"),
   704 => (x"b9",x"ff",x"49",x"bf"),
   705 => (x"66",x"c8",x"48",x"71"),
   706 => (x"58",x"a6",x"d4",x"98"),
   707 => (x"98",x"6b",x"48",x"71"),
   708 => (x"c4",x"58",x"a6",x"d0"),
   709 => (x"a6",x"c4",x"7e",x"a3"),
   710 => (x"78",x"bf",x"6e",x"48"),
   711 => (x"cc",x"48",x"66",x"d0"),
   712 => (x"c6",x"05",x"a8",x"66"),
   713 => (x"7b",x"66",x"c8",x"87"),
   714 => (x"d4",x"87",x"c6",x"c3"),
   715 => (x"ff",x"c1",x"48",x"a6"),
   716 => (x"ff",x"ff",x"ff",x"ff"),
   717 => (x"ff",x"80",x"c4",x"78"),
   718 => (x"d4",x"4a",x"c0",x"78"),
   719 => (x"49",x"72",x"4d",x"a3"),
   720 => (x"a1",x"75",x"91",x"c8"),
   721 => (x"4c",x"66",x"d0",x"49"),
   722 => (x"b7",x"c0",x"8c",x"69"),
   723 => (x"87",x"cd",x"04",x"ac"),
   724 => (x"ac",x"b7",x"66",x"d4"),
   725 => (x"dc",x"87",x"c6",x"03"),
   726 => (x"a6",x"d8",x"5a",x"a6"),
   727 => (x"c6",x"82",x"c1",x"5c"),
   728 => (x"ff",x"04",x"aa",x"b7"),
   729 => (x"66",x"d8",x"87",x"d5"),
   730 => (x"a8",x"b7",x"c0",x"48"),
   731 => (x"d8",x"87",x"d0",x"04"),
   732 => (x"91",x"c8",x"49",x"66"),
   733 => (x"21",x"49",x"a1",x"75"),
   734 => (x"69",x"48",x"6e",x"7b"),
   735 => (x"c0",x"87",x"c9",x"78"),
   736 => (x"49",x"a3",x"cc",x"7b"),
   737 => (x"78",x"69",x"48",x"6e"),
   738 => (x"6b",x"48",x"66",x"c8"),
   739 => (x"58",x"a6",x"cc",x"88"),
   740 => (x"bf",x"fc",x"ed",x"c2"),
   741 => (x"70",x"90",x"c8",x"48"),
   742 => (x"48",x"66",x"c8",x"7e"),
   743 => (x"c9",x"01",x"a8",x"6e"),
   744 => (x"48",x"66",x"c8",x"87"),
   745 => (x"c0",x"03",x"a8",x"6e"),
   746 => (x"c4",x"c1",x"87",x"fd"),
   747 => (x"bf",x"6e",x"7e",x"a3"),
   748 => (x"75",x"91",x"c8",x"49"),
   749 => (x"66",x"cc",x"49",x"a1"),
   750 => (x"49",x"bf",x"6e",x"79"),
   751 => (x"a1",x"75",x"91",x"c8"),
   752 => (x"66",x"81",x"c4",x"49"),
   753 => (x"48",x"a6",x"d0",x"79"),
   754 => (x"d0",x"78",x"bf",x"6e"),
   755 => (x"a8",x"c5",x"48",x"66"),
   756 => (x"c4",x"87",x"c7",x"05"),
   757 => (x"78",x"c0",x"48",x"a6"),
   758 => (x"66",x"d0",x"87",x"c8"),
   759 => (x"c8",x"80",x"c1",x"48"),
   760 => (x"48",x"6e",x"58",x"a6"),
   761 => (x"c8",x"78",x"66",x"c4"),
   762 => (x"49",x"73",x"1e",x"66"),
   763 => (x"c4",x"87",x"f0",x"f8"),
   764 => (x"fc",x"e5",x"c2",x"86"),
   765 => (x"f9",x"49",x"73",x"1e"),
   766 => (x"a3",x"d0",x"87",x"f2"),
   767 => (x"66",x"f0",x"c0",x"49"),
   768 => (x"26",x"8e",x"e0",x"79"),
   769 => (x"26",x"4c",x"26",x"4d"),
   770 => (x"0e",x"4f",x"26",x"4b"),
   771 => (x"0e",x"5c",x"5b",x"5e"),
   772 => (x"4b",x"c0",x"4a",x"71"),
   773 => (x"c0",x"02",x"9a",x"72"),
   774 => (x"a2",x"da",x"87",x"e0"),
   775 => (x"4b",x"69",x"9f",x"49"),
   776 => (x"bf",x"c4",x"ee",x"c2"),
   777 => (x"d4",x"87",x"cf",x"02"),
   778 => (x"69",x"9f",x"49",x"a2"),
   779 => (x"ff",x"c0",x"4c",x"49"),
   780 => (x"34",x"d0",x"9c",x"ff"),
   781 => (x"4c",x"c0",x"87",x"c2"),
   782 => (x"9b",x"73",x"b3",x"74"),
   783 => (x"4a",x"87",x"df",x"02"),
   784 => (x"ed",x"c2",x"8a",x"c2"),
   785 => (x"92",x"49",x"bf",x"fc"),
   786 => (x"bf",x"e0",x"f2",x"c2"),
   787 => (x"c2",x"80",x"72",x"48"),
   788 => (x"71",x"58",x"c0",x"f3"),
   789 => (x"c2",x"30",x"c4",x"48"),
   790 => (x"c0",x"58",x"cc",x"ee"),
   791 => (x"f2",x"c2",x"87",x"e9"),
   792 => (x"c2",x"4b",x"bf",x"e4"),
   793 => (x"c2",x"48",x"fc",x"f2"),
   794 => (x"78",x"bf",x"e8",x"f2"),
   795 => (x"bf",x"c4",x"ee",x"c2"),
   796 => (x"c2",x"87",x"c9",x"02"),
   797 => (x"49",x"bf",x"fc",x"ed"),
   798 => (x"87",x"c7",x"31",x"c4"),
   799 => (x"bf",x"ec",x"f2",x"c2"),
   800 => (x"c2",x"31",x"c4",x"49"),
   801 => (x"c2",x"59",x"cc",x"ee"),
   802 => (x"26",x"5b",x"fc",x"f2"),
   803 => (x"26",x"4b",x"26",x"4c"),
   804 => (x"5b",x"5e",x"0e",x"4f"),
   805 => (x"f0",x"0e",x"5d",x"5c"),
   806 => (x"59",x"a6",x"c8",x"86"),
   807 => (x"ff",x"ff",x"ff",x"cf"),
   808 => (x"7e",x"c0",x"4c",x"f8"),
   809 => (x"d8",x"02",x"66",x"c4"),
   810 => (x"f8",x"e5",x"c2",x"87"),
   811 => (x"c2",x"78",x"c0",x"48"),
   812 => (x"c2",x"48",x"f0",x"e5"),
   813 => (x"78",x"bf",x"fc",x"f2"),
   814 => (x"48",x"f4",x"e5",x"c2"),
   815 => (x"bf",x"f8",x"f2",x"c2"),
   816 => (x"d9",x"ee",x"c2",x"78"),
   817 => (x"c2",x"50",x"c0",x"48"),
   818 => (x"49",x"bf",x"c8",x"ee"),
   819 => (x"bf",x"f8",x"e5",x"c2"),
   820 => (x"03",x"aa",x"71",x"4a"),
   821 => (x"72",x"87",x"cc",x"c4"),
   822 => (x"05",x"99",x"cf",x"49"),
   823 => (x"c0",x"87",x"ea",x"c0"),
   824 => (x"c2",x"48",x"cc",x"fa"),
   825 => (x"78",x"bf",x"f0",x"e5"),
   826 => (x"1e",x"fc",x"e5",x"c2"),
   827 => (x"bf",x"f0",x"e5",x"c2"),
   828 => (x"f0",x"e5",x"c2",x"49"),
   829 => (x"78",x"a1",x"c1",x"48"),
   830 => (x"f9",x"df",x"ff",x"71"),
   831 => (x"c0",x"86",x"c4",x"87"),
   832 => (x"c2",x"48",x"c8",x"fa"),
   833 => (x"cc",x"78",x"fc",x"e5"),
   834 => (x"c8",x"fa",x"c0",x"87"),
   835 => (x"e0",x"c0",x"48",x"bf"),
   836 => (x"cc",x"fa",x"c0",x"80"),
   837 => (x"f8",x"e5",x"c2",x"58"),
   838 => (x"80",x"c1",x"48",x"bf"),
   839 => (x"58",x"fc",x"e5",x"c2"),
   840 => (x"00",x"0e",x"88",x"27"),
   841 => (x"bf",x"97",x"bf",x"00"),
   842 => (x"c2",x"02",x"9d",x"4d"),
   843 => (x"e5",x"c3",x"87",x"e5"),
   844 => (x"de",x"c2",x"02",x"ad"),
   845 => (x"c8",x"fa",x"c0",x"87"),
   846 => (x"a3",x"cb",x"4b",x"bf"),
   847 => (x"cf",x"4c",x"11",x"49"),
   848 => (x"d2",x"c1",x"05",x"ac"),
   849 => (x"df",x"49",x"75",x"87"),
   850 => (x"cd",x"89",x"c1",x"99"),
   851 => (x"cc",x"ee",x"c2",x"91"),
   852 => (x"4a",x"a3",x"c1",x"81"),
   853 => (x"a3",x"c3",x"51",x"12"),
   854 => (x"c5",x"51",x"12",x"4a"),
   855 => (x"51",x"12",x"4a",x"a3"),
   856 => (x"12",x"4a",x"a3",x"c7"),
   857 => (x"4a",x"a3",x"c9",x"51"),
   858 => (x"a3",x"ce",x"51",x"12"),
   859 => (x"d0",x"51",x"12",x"4a"),
   860 => (x"51",x"12",x"4a",x"a3"),
   861 => (x"12",x"4a",x"a3",x"d2"),
   862 => (x"4a",x"a3",x"d4",x"51"),
   863 => (x"a3",x"d6",x"51",x"12"),
   864 => (x"d8",x"51",x"12",x"4a"),
   865 => (x"51",x"12",x"4a",x"a3"),
   866 => (x"12",x"4a",x"a3",x"dc"),
   867 => (x"4a",x"a3",x"de",x"51"),
   868 => (x"7e",x"c1",x"51",x"12"),
   869 => (x"74",x"87",x"fc",x"c0"),
   870 => (x"05",x"99",x"c8",x"49"),
   871 => (x"74",x"87",x"ed",x"c0"),
   872 => (x"05",x"99",x"d0",x"49"),
   873 => (x"e0",x"c0",x"87",x"d3"),
   874 => (x"cc",x"c0",x"02",x"66"),
   875 => (x"c0",x"49",x"73",x"87"),
   876 => (x"70",x"0f",x"66",x"e0"),
   877 => (x"d3",x"c0",x"02",x"98"),
   878 => (x"c0",x"05",x"6e",x"87"),
   879 => (x"ee",x"c2",x"87",x"c6"),
   880 => (x"50",x"c0",x"48",x"cc"),
   881 => (x"bf",x"c8",x"fa",x"c0"),
   882 => (x"87",x"e9",x"c2",x"48"),
   883 => (x"48",x"d9",x"ee",x"c2"),
   884 => (x"c2",x"7e",x"50",x"c0"),
   885 => (x"49",x"bf",x"c8",x"ee"),
   886 => (x"bf",x"f8",x"e5",x"c2"),
   887 => (x"04",x"aa",x"71",x"4a"),
   888 => (x"cf",x"87",x"f4",x"fb"),
   889 => (x"f8",x"ff",x"ff",x"ff"),
   890 => (x"fc",x"f2",x"c2",x"4c"),
   891 => (x"c8",x"c0",x"05",x"bf"),
   892 => (x"c4",x"ee",x"c2",x"87"),
   893 => (x"fa",x"c1",x"02",x"bf"),
   894 => (x"f4",x"e5",x"c2",x"87"),
   895 => (x"c0",x"eb",x"49",x"bf"),
   896 => (x"f8",x"e5",x"c2",x"87"),
   897 => (x"48",x"a6",x"c4",x"58"),
   898 => (x"bf",x"f4",x"e5",x"c2"),
   899 => (x"c4",x"ee",x"c2",x"78"),
   900 => (x"db",x"c0",x"02",x"bf"),
   901 => (x"49",x"66",x"c4",x"87"),
   902 => (x"a9",x"74",x"99",x"74"),
   903 => (x"87",x"c8",x"c0",x"02"),
   904 => (x"c0",x"48",x"a6",x"c8"),
   905 => (x"87",x"e7",x"c0",x"78"),
   906 => (x"c1",x"48",x"a6",x"c8"),
   907 => (x"87",x"df",x"c0",x"78"),
   908 => (x"cf",x"49",x"66",x"c4"),
   909 => (x"a9",x"99",x"f8",x"ff"),
   910 => (x"87",x"c8",x"c0",x"02"),
   911 => (x"c0",x"48",x"a6",x"cc"),
   912 => (x"87",x"c5",x"c0",x"78"),
   913 => (x"c1",x"48",x"a6",x"cc"),
   914 => (x"48",x"a6",x"c8",x"78"),
   915 => (x"c8",x"78",x"66",x"cc"),
   916 => (x"de",x"c0",x"05",x"66"),
   917 => (x"49",x"66",x"c4",x"87"),
   918 => (x"ed",x"c2",x"89",x"c2"),
   919 => (x"c2",x"91",x"bf",x"fc"),
   920 => (x"48",x"bf",x"e0",x"f2"),
   921 => (x"e5",x"c2",x"80",x"71"),
   922 => (x"e5",x"c2",x"58",x"f4"),
   923 => (x"78",x"c0",x"48",x"f8"),
   924 => (x"c0",x"87",x"d4",x"f9"),
   925 => (x"ff",x"ff",x"cf",x"48"),
   926 => (x"f0",x"4c",x"f8",x"ff"),
   927 => (x"26",x"4d",x"26",x"8e"),
   928 => (x"26",x"4b",x"26",x"4c"),
   929 => (x"00",x"00",x"00",x"4f"),
   930 => (x"00",x"00",x"00",x"00"),
   931 => (x"ff",x"ff",x"ff",x"ff"),
   932 => (x"48",x"d4",x"ff",x"1e"),
   933 => (x"68",x"78",x"ff",x"c3"),
   934 => (x"1e",x"4f",x"26",x"48"),
   935 => (x"c3",x"48",x"d4",x"ff"),
   936 => (x"d0",x"ff",x"78",x"ff"),
   937 => (x"78",x"e1",x"c0",x"48"),
   938 => (x"d4",x"48",x"d4",x"ff"),
   939 => (x"1e",x"4f",x"26",x"78"),
   940 => (x"c0",x"48",x"d0",x"ff"),
   941 => (x"4f",x"26",x"78",x"e0"),
   942 => (x"87",x"d4",x"ff",x"1e"),
   943 => (x"02",x"99",x"49",x"70"),
   944 => (x"fb",x"c0",x"87",x"c6"),
   945 => (x"87",x"f1",x"05",x"a9"),
   946 => (x"4f",x"26",x"48",x"71"),
   947 => (x"5c",x"5b",x"5e",x"0e"),
   948 => (x"c0",x"4b",x"71",x"0e"),
   949 => (x"87",x"f8",x"fe",x"4c"),
   950 => (x"02",x"99",x"49",x"70"),
   951 => (x"c0",x"87",x"f9",x"c0"),
   952 => (x"c0",x"02",x"a9",x"ec"),
   953 => (x"fb",x"c0",x"87",x"f2"),
   954 => (x"eb",x"c0",x"02",x"a9"),
   955 => (x"b7",x"66",x"cc",x"87"),
   956 => (x"87",x"c7",x"03",x"ac"),
   957 => (x"c2",x"02",x"66",x"d0"),
   958 => (x"71",x"53",x"71",x"87"),
   959 => (x"87",x"c2",x"02",x"99"),
   960 => (x"cb",x"fe",x"84",x"c1"),
   961 => (x"99",x"49",x"70",x"87"),
   962 => (x"c0",x"87",x"cd",x"02"),
   963 => (x"c7",x"02",x"a9",x"ec"),
   964 => (x"a9",x"fb",x"c0",x"87"),
   965 => (x"87",x"d5",x"ff",x"05"),
   966 => (x"c3",x"02",x"66",x"d0"),
   967 => (x"7b",x"97",x"c0",x"87"),
   968 => (x"05",x"a9",x"ec",x"c0"),
   969 => (x"4a",x"74",x"87",x"c4"),
   970 => (x"4a",x"74",x"87",x"c5"),
   971 => (x"72",x"8a",x"0a",x"c0"),
   972 => (x"26",x"4c",x"26",x"48"),
   973 => (x"1e",x"4f",x"26",x"4b"),
   974 => (x"70",x"87",x"d5",x"fd"),
   975 => (x"a9",x"f0",x"c0",x"49"),
   976 => (x"c0",x"87",x"c9",x"04"),
   977 => (x"c3",x"01",x"a9",x"f9"),
   978 => (x"89",x"f0",x"c0",x"87"),
   979 => (x"04",x"a9",x"c1",x"c1"),
   980 => (x"da",x"c1",x"87",x"c9"),
   981 => (x"87",x"c3",x"01",x"a9"),
   982 => (x"71",x"89",x"f7",x"c0"),
   983 => (x"0e",x"4f",x"26",x"48"),
   984 => (x"5d",x"5c",x"5b",x"5e"),
   985 => (x"71",x"86",x"f8",x"0e"),
   986 => (x"fc",x"7e",x"c0",x"4c"),
   987 => (x"4b",x"c0",x"87",x"ed"),
   988 => (x"97",x"c0",x"c0",x"c1"),
   989 => (x"a9",x"c0",x"49",x"bf"),
   990 => (x"fc",x"87",x"cf",x"04"),
   991 => (x"83",x"c1",x"87",x"fa"),
   992 => (x"97",x"c0",x"c0",x"c1"),
   993 => (x"06",x"ab",x"49",x"bf"),
   994 => (x"c0",x"c1",x"87",x"f1"),
   995 => (x"02",x"bf",x"97",x"c0"),
   996 => (x"fb",x"fb",x"87",x"cf"),
   997 => (x"99",x"49",x"70",x"87"),
   998 => (x"c0",x"87",x"c6",x"02"),
   999 => (x"f1",x"05",x"a9",x"ec"),
  1000 => (x"fb",x"4b",x"c0",x"87"),
  1001 => (x"4d",x"70",x"87",x"ea"),
  1002 => (x"c8",x"87",x"e5",x"fb"),
  1003 => (x"df",x"fb",x"58",x"a6"),
  1004 => (x"c1",x"4a",x"70",x"87"),
  1005 => (x"49",x"a4",x"c8",x"83"),
  1006 => (x"ad",x"49",x"69",x"97"),
  1007 => (x"c9",x"87",x"da",x"05"),
  1008 => (x"69",x"97",x"49",x"a4"),
  1009 => (x"a9",x"66",x"c4",x"49"),
  1010 => (x"ca",x"87",x"ce",x"05"),
  1011 => (x"69",x"97",x"49",x"a4"),
  1012 => (x"c4",x"05",x"aa",x"49"),
  1013 => (x"d0",x"7e",x"c1",x"87"),
  1014 => (x"ad",x"ec",x"c0",x"87"),
  1015 => (x"c0",x"87",x"c6",x"02"),
  1016 => (x"c4",x"05",x"ad",x"fb"),
  1017 => (x"c1",x"4b",x"c0",x"87"),
  1018 => (x"fe",x"02",x"6e",x"7e"),
  1019 => (x"fe",x"fa",x"87",x"f5"),
  1020 => (x"f8",x"48",x"73",x"87"),
  1021 => (x"26",x"4d",x"26",x"8e"),
  1022 => (x"26",x"4b",x"26",x"4c"),
  1023 => (x"00",x"00",x"00",x"4f"),
  1024 => (x"1e",x"73",x"1e",x"00"),
  1025 => (x"c8",x"4b",x"d4",x"ff"),
  1026 => (x"d0",x"ff",x"4a",x"66"),
  1027 => (x"78",x"c5",x"c8",x"48"),
  1028 => (x"c1",x"48",x"d4",x"ff"),
  1029 => (x"7b",x"11",x"78",x"d4"),
  1030 => (x"f9",x"05",x"8a",x"c1"),
  1031 => (x"48",x"d0",x"ff",x"87"),
  1032 => (x"4b",x"26",x"78",x"c4"),
  1033 => (x"5e",x"0e",x"4f",x"26"),
  1034 => (x"0e",x"5d",x"5c",x"5b"),
  1035 => (x"7e",x"71",x"86",x"f8"),
  1036 => (x"f3",x"c2",x"1e",x"6e"),
  1037 => (x"ff",x"e3",x"49",x"d0"),
  1038 => (x"70",x"86",x"c4",x"87"),
  1039 => (x"e4",x"c4",x"02",x"98"),
  1040 => (x"e8",x"ed",x"c1",x"87"),
  1041 => (x"49",x"6e",x"4c",x"bf"),
  1042 => (x"c8",x"87",x"d4",x"fc"),
  1043 => (x"98",x"70",x"58",x"a6"),
  1044 => (x"c4",x"87",x"c5",x"05"),
  1045 => (x"78",x"c1",x"48",x"a6"),
  1046 => (x"c5",x"48",x"d0",x"ff"),
  1047 => (x"48",x"d4",x"ff",x"78"),
  1048 => (x"c4",x"78",x"d5",x"c1"),
  1049 => (x"89",x"c1",x"49",x"66"),
  1050 => (x"ed",x"c1",x"31",x"c6"),
  1051 => (x"4a",x"bf",x"97",x"e0"),
  1052 => (x"ff",x"b0",x"71",x"48"),
  1053 => (x"ff",x"78",x"08",x"d4"),
  1054 => (x"78",x"c4",x"48",x"d0"),
  1055 => (x"97",x"cc",x"f3",x"c2"),
  1056 => (x"99",x"d0",x"49",x"bf"),
  1057 => (x"c5",x"87",x"dd",x"02"),
  1058 => (x"48",x"d4",x"ff",x"78"),
  1059 => (x"c0",x"78",x"d6",x"c1"),
  1060 => (x"48",x"d4",x"ff",x"4a"),
  1061 => (x"c1",x"78",x"ff",x"c3"),
  1062 => (x"aa",x"e0",x"c0",x"82"),
  1063 => (x"ff",x"87",x"f2",x"04"),
  1064 => (x"78",x"c4",x"48",x"d0"),
  1065 => (x"c3",x"48",x"d4",x"ff"),
  1066 => (x"d0",x"ff",x"78",x"ff"),
  1067 => (x"ff",x"78",x"c5",x"48"),
  1068 => (x"d3",x"c1",x"48",x"d4"),
  1069 => (x"ff",x"78",x"c1",x"78"),
  1070 => (x"78",x"c4",x"48",x"d0"),
  1071 => (x"06",x"ac",x"b7",x"c0"),
  1072 => (x"c2",x"87",x"cb",x"c2"),
  1073 => (x"4b",x"bf",x"d8",x"f3"),
  1074 => (x"73",x"7e",x"74",x"8c"),
  1075 => (x"dd",x"c1",x"02",x"9b"),
  1076 => (x"4d",x"c0",x"c8",x"87"),
  1077 => (x"ab",x"b7",x"c0",x"8b"),
  1078 => (x"c8",x"87",x"c6",x"03"),
  1079 => (x"c0",x"4d",x"a3",x"c0"),
  1080 => (x"cc",x"f3",x"c2",x"4b"),
  1081 => (x"d0",x"49",x"bf",x"97"),
  1082 => (x"87",x"cf",x"02",x"99"),
  1083 => (x"f3",x"c2",x"1e",x"c0"),
  1084 => (x"f7",x"e5",x"49",x"d0"),
  1085 => (x"70",x"86",x"c4",x"87"),
  1086 => (x"c2",x"87",x"d8",x"4c"),
  1087 => (x"c2",x"1e",x"fc",x"e5"),
  1088 => (x"e5",x"49",x"d0",x"f3"),
  1089 => (x"4c",x"70",x"87",x"e6"),
  1090 => (x"e5",x"c2",x"1e",x"75"),
  1091 => (x"f0",x"fb",x"49",x"fc"),
  1092 => (x"74",x"86",x"c8",x"87"),
  1093 => (x"87",x"c5",x"05",x"9c"),
  1094 => (x"ca",x"c1",x"48",x"c0"),
  1095 => (x"c2",x"1e",x"c1",x"87"),
  1096 => (x"e3",x"49",x"d0",x"f3"),
  1097 => (x"86",x"c4",x"87",x"f9"),
  1098 => (x"fe",x"05",x"9b",x"73"),
  1099 => (x"4c",x"6e",x"87",x"e3"),
  1100 => (x"06",x"ac",x"b7",x"c0"),
  1101 => (x"f3",x"c2",x"87",x"d1"),
  1102 => (x"78",x"c0",x"48",x"d0"),
  1103 => (x"78",x"c0",x"80",x"d0"),
  1104 => (x"f3",x"c2",x"80",x"f4"),
  1105 => (x"c0",x"78",x"bf",x"dc"),
  1106 => (x"fd",x"01",x"ac",x"b7"),
  1107 => (x"d0",x"ff",x"87",x"f5"),
  1108 => (x"ff",x"78",x"c5",x"48"),
  1109 => (x"d3",x"c1",x"48",x"d4"),
  1110 => (x"ff",x"78",x"c0",x"78"),
  1111 => (x"78",x"c4",x"48",x"d0"),
  1112 => (x"c2",x"c0",x"48",x"c1"),
  1113 => (x"f8",x"48",x"c0",x"87"),
  1114 => (x"26",x"4d",x"26",x"8e"),
  1115 => (x"26",x"4b",x"26",x"4c"),
  1116 => (x"5b",x"5e",x"0e",x"4f"),
  1117 => (x"fc",x"0e",x"5d",x"5c"),
  1118 => (x"c0",x"4d",x"71",x"86"),
  1119 => (x"04",x"ad",x"4c",x"4b"),
  1120 => (x"c0",x"87",x"e8",x"c0"),
  1121 => (x"74",x"1e",x"df",x"fd"),
  1122 => (x"87",x"c4",x"02",x"9c"),
  1123 => (x"87",x"c2",x"4a",x"c0"),
  1124 => (x"49",x"72",x"4a",x"c1"),
  1125 => (x"c4",x"87",x"fa",x"eb"),
  1126 => (x"c1",x"7e",x"70",x"86"),
  1127 => (x"c2",x"05",x"6e",x"83"),
  1128 => (x"c1",x"4b",x"75",x"87"),
  1129 => (x"06",x"ab",x"75",x"84"),
  1130 => (x"6e",x"87",x"d8",x"ff"),
  1131 => (x"26",x"8e",x"fc",x"48"),
  1132 => (x"26",x"4c",x"26",x"4d"),
  1133 => (x"0e",x"4f",x"26",x"4b"),
  1134 => (x"0e",x"5c",x"5b",x"5e"),
  1135 => (x"66",x"cc",x"4b",x"71"),
  1136 => (x"4c",x"87",x"d8",x"02"),
  1137 => (x"02",x"8c",x"f0",x"c0"),
  1138 => (x"4a",x"74",x"87",x"d8"),
  1139 => (x"d1",x"02",x"8a",x"c1"),
  1140 => (x"cd",x"02",x"8a",x"87"),
  1141 => (x"c9",x"02",x"8a",x"87"),
  1142 => (x"73",x"87",x"d9",x"87"),
  1143 => (x"87",x"c6",x"f9",x"49"),
  1144 => (x"1e",x"74",x"87",x"d2"),
  1145 => (x"da",x"c1",x"49",x"c0"),
  1146 => (x"1e",x"74",x"87",x"f6"),
  1147 => (x"da",x"c1",x"49",x"73"),
  1148 => (x"86",x"c8",x"87",x"ee"),
  1149 => (x"4b",x"26",x"4c",x"26"),
  1150 => (x"5e",x"0e",x"4f",x"26"),
  1151 => (x"0e",x"5d",x"5c",x"5b"),
  1152 => (x"4c",x"71",x"86",x"fc"),
  1153 => (x"c2",x"91",x"de",x"49"),
  1154 => (x"71",x"4d",x"f0",x"f4"),
  1155 => (x"02",x"6d",x"97",x"85"),
  1156 => (x"c2",x"87",x"dc",x"c1"),
  1157 => (x"49",x"bf",x"e0",x"f4"),
  1158 => (x"fd",x"71",x"81",x"74"),
  1159 => (x"7e",x"70",x"87",x"d3"),
  1160 => (x"c0",x"02",x"98",x"48"),
  1161 => (x"f4",x"c2",x"87",x"f2"),
  1162 => (x"4a",x"70",x"4b",x"e4"),
  1163 => (x"fb",x"fe",x"49",x"cb"),
  1164 => (x"4b",x"74",x"87",x"f1"),
  1165 => (x"ed",x"c1",x"93",x"cc"),
  1166 => (x"83",x"c4",x"83",x"ec"),
  1167 => (x"7b",x"fc",x"c9",x"c1"),
  1168 => (x"c2",x"c1",x"49",x"74"),
  1169 => (x"7b",x"75",x"87",x"fa"),
  1170 => (x"97",x"e4",x"ed",x"c1"),
  1171 => (x"c2",x"1e",x"49",x"bf"),
  1172 => (x"fd",x"49",x"e4",x"f4"),
  1173 => (x"86",x"c4",x"87",x"e1"),
  1174 => (x"c2",x"c1",x"49",x"74"),
  1175 => (x"49",x"c0",x"87",x"e2"),
  1176 => (x"87",x"fd",x"c3",x"c1"),
  1177 => (x"48",x"c8",x"f3",x"c2"),
  1178 => (x"c0",x"49",x"50",x"c0"),
  1179 => (x"fc",x"87",x"c3",x"e1"),
  1180 => (x"26",x"4d",x"26",x"8e"),
  1181 => (x"26",x"4b",x"26",x"4c"),
  1182 => (x"00",x"00",x"00",x"4f"),
  1183 => (x"64",x"61",x"6f",x"4c"),
  1184 => (x"2e",x"67",x"6e",x"69"),
  1185 => (x"00",x"00",x"2e",x"2e"),
  1186 => (x"61",x"42",x"20",x"80"),
  1187 => (x"00",x"00",x"6b",x"63"),
  1188 => (x"64",x"61",x"6f",x"4c"),
  1189 => (x"20",x"2e",x"2a",x"20"),
  1190 => (x"00",x"00",x"00",x"00"),
  1191 => (x"00",x"00",x"20",x"3a"),
  1192 => (x"61",x"42",x"20",x"80"),
  1193 => (x"00",x"00",x"6b",x"63"),
  1194 => (x"78",x"45",x"20",x"80"),
  1195 => (x"00",x"00",x"74",x"69"),
  1196 => (x"49",x"20",x"44",x"53"),
  1197 => (x"2e",x"74",x"69",x"6e"),
  1198 => (x"00",x"00",x"00",x"2e"),
  1199 => (x"00",x"00",x"4b",x"4f"),
  1200 => (x"54",x"4f",x"4f",x"42"),
  1201 => (x"20",x"20",x"20",x"20"),
  1202 => (x"00",x"4d",x"4f",x"52"),
  1203 => (x"71",x"1e",x"73",x"1e"),
  1204 => (x"f4",x"c2",x"49",x"4b"),
  1205 => (x"71",x"81",x"bf",x"e0"),
  1206 => (x"70",x"87",x"d6",x"fa"),
  1207 => (x"c4",x"02",x"9a",x"4a"),
  1208 => (x"e6",x"e4",x"49",x"87"),
  1209 => (x"e0",x"f4",x"c2",x"87"),
  1210 => (x"73",x"78",x"c0",x"48"),
  1211 => (x"87",x"fa",x"c1",x"49"),
  1212 => (x"4f",x"26",x"4b",x"26"),
  1213 => (x"71",x"1e",x"73",x"1e"),
  1214 => (x"4a",x"a3",x"c4",x"4b"),
  1215 => (x"87",x"d0",x"c1",x"02"),
  1216 => (x"dc",x"02",x"8a",x"c1"),
  1217 => (x"c0",x"02",x"8a",x"87"),
  1218 => (x"05",x"8a",x"87",x"f2"),
  1219 => (x"c2",x"87",x"d3",x"c1"),
  1220 => (x"02",x"bf",x"e0",x"f4"),
  1221 => (x"48",x"87",x"cb",x"c1"),
  1222 => (x"f4",x"c2",x"88",x"c1"),
  1223 => (x"c1",x"c1",x"58",x"e4"),
  1224 => (x"e0",x"f4",x"c2",x"87"),
  1225 => (x"89",x"c6",x"49",x"bf"),
  1226 => (x"59",x"e4",x"f4",x"c2"),
  1227 => (x"03",x"a9",x"b7",x"c0"),
  1228 => (x"c2",x"87",x"ef",x"c0"),
  1229 => (x"c0",x"48",x"e0",x"f4"),
  1230 => (x"87",x"e6",x"c0",x"78"),
  1231 => (x"bf",x"dc",x"f4",x"c2"),
  1232 => (x"c2",x"87",x"df",x"02"),
  1233 => (x"48",x"bf",x"e0",x"f4"),
  1234 => (x"f4",x"c2",x"80",x"c1"),
  1235 => (x"87",x"d2",x"58",x"e4"),
  1236 => (x"bf",x"dc",x"f4",x"c2"),
  1237 => (x"c2",x"87",x"cb",x"02"),
  1238 => (x"48",x"bf",x"e0",x"f4"),
  1239 => (x"f4",x"c2",x"80",x"c6"),
  1240 => (x"49",x"73",x"58",x"e4"),
  1241 => (x"4b",x"26",x"87",x"c4"),
  1242 => (x"5e",x"0e",x"4f",x"26"),
  1243 => (x"0e",x"5d",x"5c",x"5b"),
  1244 => (x"a6",x"d0",x"86",x"f0"),
  1245 => (x"fc",x"e5",x"c2",x"59"),
  1246 => (x"c2",x"4c",x"c0",x"4d"),
  1247 => (x"c1",x"48",x"dc",x"f4"),
  1248 => (x"48",x"a6",x"c8",x"78"),
  1249 => (x"7e",x"75",x"78",x"c0"),
  1250 => (x"bf",x"e0",x"f4",x"c2"),
  1251 => (x"06",x"a8",x"c0",x"48"),
  1252 => (x"c8",x"87",x"c0",x"c1"),
  1253 => (x"7e",x"75",x"5c",x"a6"),
  1254 => (x"48",x"fc",x"e5",x"c2"),
  1255 => (x"f2",x"c0",x"02",x"98"),
  1256 => (x"4d",x"66",x"c4",x"87"),
  1257 => (x"1e",x"df",x"fd",x"c0"),
  1258 => (x"c4",x"02",x"66",x"cc"),
  1259 => (x"c2",x"4c",x"c0",x"87"),
  1260 => (x"74",x"4c",x"c1",x"87"),
  1261 => (x"87",x"d9",x"e3",x"49"),
  1262 => (x"7e",x"70",x"86",x"c4"),
  1263 => (x"66",x"c8",x"85",x"c1"),
  1264 => (x"cc",x"80",x"c1",x"48"),
  1265 => (x"f4",x"c2",x"58",x"a6"),
  1266 => (x"03",x"ad",x"bf",x"e0"),
  1267 => (x"05",x"6e",x"87",x"c5"),
  1268 => (x"6e",x"87",x"d1",x"ff"),
  1269 => (x"75",x"4c",x"c0",x"4d"),
  1270 => (x"dc",x"c3",x"02",x"9d"),
  1271 => (x"df",x"fd",x"c0",x"87"),
  1272 => (x"02",x"66",x"cc",x"1e"),
  1273 => (x"a6",x"c8",x"87",x"c7"),
  1274 => (x"c5",x"78",x"c0",x"48"),
  1275 => (x"48",x"a6",x"c8",x"87"),
  1276 => (x"66",x"c8",x"78",x"c1"),
  1277 => (x"87",x"d9",x"e2",x"49"),
  1278 => (x"7e",x"70",x"86",x"c4"),
  1279 => (x"c2",x"02",x"98",x"48"),
  1280 => (x"cb",x"49",x"87",x"e4"),
  1281 => (x"49",x"69",x"97",x"81"),
  1282 => (x"c1",x"02",x"99",x"d0"),
  1283 => (x"49",x"74",x"87",x"d4"),
  1284 => (x"ed",x"c1",x"91",x"cc"),
  1285 => (x"cb",x"c1",x"81",x"ec"),
  1286 => (x"81",x"c8",x"79",x"cc"),
  1287 => (x"74",x"51",x"ff",x"c3"),
  1288 => (x"c2",x"91",x"de",x"49"),
  1289 => (x"71",x"4d",x"f0",x"f4"),
  1290 => (x"97",x"c1",x"c2",x"85"),
  1291 => (x"49",x"a5",x"c1",x"7d"),
  1292 => (x"c2",x"51",x"e0",x"c0"),
  1293 => (x"bf",x"97",x"cc",x"ee"),
  1294 => (x"c1",x"87",x"d2",x"02"),
  1295 => (x"4b",x"a5",x"c2",x"84"),
  1296 => (x"4a",x"cc",x"ee",x"c2"),
  1297 => (x"f3",x"fe",x"49",x"db"),
  1298 => (x"d9",x"c1",x"87",x"d9"),
  1299 => (x"49",x"a5",x"cd",x"87"),
  1300 => (x"84",x"c1",x"51",x"c0"),
  1301 => (x"6e",x"4b",x"a5",x"c2"),
  1302 => (x"fe",x"49",x"cb",x"4a"),
  1303 => (x"c1",x"87",x"c4",x"f3"),
  1304 => (x"49",x"74",x"87",x"c4"),
  1305 => (x"ed",x"c1",x"91",x"cc"),
  1306 => (x"c7",x"c1",x"81",x"ec"),
  1307 => (x"ee",x"c2",x"79",x"fa"),
  1308 => (x"02",x"bf",x"97",x"cc"),
  1309 => (x"49",x"74",x"87",x"d8"),
  1310 => (x"84",x"c1",x"91",x"de"),
  1311 => (x"4b",x"f0",x"f4",x"c2"),
  1312 => (x"ee",x"c2",x"83",x"71"),
  1313 => (x"49",x"dd",x"4a",x"cc"),
  1314 => (x"87",x"d7",x"f2",x"fe"),
  1315 => (x"4b",x"74",x"87",x"d8"),
  1316 => (x"f4",x"c2",x"93",x"de"),
  1317 => (x"a3",x"cb",x"83",x"f0"),
  1318 => (x"c1",x"51",x"c0",x"49"),
  1319 => (x"4a",x"6e",x"73",x"84"),
  1320 => (x"f1",x"fe",x"49",x"cb"),
  1321 => (x"66",x"c8",x"87",x"fd"),
  1322 => (x"cc",x"80",x"c1",x"48"),
  1323 => (x"ac",x"c7",x"58",x"a6"),
  1324 => (x"87",x"c5",x"c0",x"03"),
  1325 => (x"e4",x"fc",x"05",x"6e"),
  1326 => (x"03",x"ac",x"c7",x"87"),
  1327 => (x"c2",x"87",x"e4",x"c0"),
  1328 => (x"c0",x"48",x"dc",x"f4"),
  1329 => (x"cc",x"49",x"74",x"78"),
  1330 => (x"ec",x"ed",x"c1",x"91"),
  1331 => (x"fa",x"c7",x"c1",x"81"),
  1332 => (x"de",x"49",x"74",x"79"),
  1333 => (x"f0",x"f4",x"c2",x"91"),
  1334 => (x"c1",x"51",x"c0",x"81"),
  1335 => (x"04",x"ac",x"c7",x"84"),
  1336 => (x"c1",x"87",x"dc",x"ff"),
  1337 => (x"c0",x"48",x"c8",x"ef"),
  1338 => (x"c1",x"80",x"f7",x"50"),
  1339 => (x"c1",x"40",x"d0",x"d5"),
  1340 => (x"c8",x"78",x"c8",x"ca"),
  1341 => (x"f4",x"cb",x"c1",x"80"),
  1342 => (x"49",x"66",x"cc",x"78"),
  1343 => (x"87",x"c0",x"f8",x"c0"),
  1344 => (x"4d",x"26",x"8e",x"f0"),
  1345 => (x"4b",x"26",x"4c",x"26"),
  1346 => (x"73",x"1e",x"4f",x"26"),
  1347 => (x"49",x"4b",x"71",x"1e"),
  1348 => (x"ed",x"c1",x"91",x"cc"),
  1349 => (x"a1",x"c8",x"81",x"ec"),
  1350 => (x"e0",x"ed",x"c1",x"4a"),
  1351 => (x"c9",x"50",x"12",x"48"),
  1352 => (x"c0",x"c1",x"4a",x"a1"),
  1353 => (x"50",x"12",x"48",x"c0"),
  1354 => (x"ed",x"c1",x"81",x"ca"),
  1355 => (x"50",x"11",x"48",x"e4"),
  1356 => (x"97",x"e4",x"ed",x"c1"),
  1357 => (x"c0",x"1e",x"49",x"bf"),
  1358 => (x"87",x"fb",x"f1",x"49"),
  1359 => (x"e9",x"f8",x"49",x"73"),
  1360 => (x"26",x"8e",x"fc",x"87"),
  1361 => (x"1e",x"4f",x"26",x"4b"),
  1362 => (x"f8",x"c0",x"49",x"c0"),
  1363 => (x"4f",x"26",x"87",x"d3"),
  1364 => (x"49",x"4a",x"71",x"1e"),
  1365 => (x"ed",x"c1",x"91",x"cc"),
  1366 => (x"81",x"c8",x"81",x"ec"),
  1367 => (x"48",x"c8",x"f3",x"c2"),
  1368 => (x"f0",x"c0",x"50",x"11"),
  1369 => (x"ec",x"fe",x"49",x"a2"),
  1370 => (x"49",x"c0",x"87",x"e2"),
  1371 => (x"26",x"87",x"c3",x"d5"),
  1372 => (x"d4",x"ff",x"1e",x"4f"),
  1373 => (x"7a",x"ff",x"c3",x"4a"),
  1374 => (x"c0",x"48",x"d0",x"ff"),
  1375 => (x"7a",x"de",x"78",x"e1"),
  1376 => (x"c8",x"48",x"7a",x"71"),
  1377 => (x"7a",x"70",x"28",x"b7"),
  1378 => (x"b7",x"d0",x"48",x"71"),
  1379 => (x"71",x"7a",x"70",x"28"),
  1380 => (x"28",x"b7",x"d8",x"48"),
  1381 => (x"d0",x"ff",x"7a",x"70"),
  1382 => (x"78",x"e0",x"c0",x"48"),
  1383 => (x"5e",x"0e",x"4f",x"26"),
  1384 => (x"0e",x"5d",x"5c",x"5b"),
  1385 => (x"4d",x"71",x"86",x"f4"),
  1386 => (x"c1",x"91",x"cc",x"49"),
  1387 => (x"c8",x"81",x"ec",x"ed"),
  1388 => (x"a1",x"ca",x"4a",x"a1"),
  1389 => (x"48",x"a6",x"c4",x"7e"),
  1390 => (x"bf",x"c4",x"f3",x"c2"),
  1391 => (x"bf",x"97",x"6e",x"78"),
  1392 => (x"4c",x"66",x"c4",x"4b"),
  1393 => (x"48",x"12",x"2c",x"73"),
  1394 => (x"70",x"58",x"a6",x"cc"),
  1395 => (x"c9",x"84",x"c1",x"9c"),
  1396 => (x"49",x"69",x"97",x"81"),
  1397 => (x"c2",x"04",x"ac",x"b7"),
  1398 => (x"6e",x"4c",x"c0",x"87"),
  1399 => (x"c8",x"4a",x"bf",x"97"),
  1400 => (x"31",x"72",x"49",x"66"),
  1401 => (x"66",x"c4",x"b9",x"ff"),
  1402 => (x"72",x"48",x"74",x"99"),
  1403 => (x"b1",x"4a",x"70",x"30"),
  1404 => (x"59",x"c8",x"f3",x"c2"),
  1405 => (x"87",x"f9",x"fd",x"71"),
  1406 => (x"f4",x"c2",x"1e",x"c7"),
  1407 => (x"c1",x"1e",x"bf",x"d8"),
  1408 => (x"c2",x"1e",x"ec",x"ed"),
  1409 => (x"bf",x"97",x"c8",x"f3"),
  1410 => (x"87",x"f4",x"c1",x"49"),
  1411 => (x"f3",x"c0",x"49",x"75"),
  1412 => (x"8e",x"e8",x"87",x"ee"),
  1413 => (x"4c",x"26",x"4d",x"26"),
  1414 => (x"4f",x"26",x"4b",x"26"),
  1415 => (x"71",x"1e",x"73",x"1e"),
  1416 => (x"f9",x"fd",x"49",x"4b"),
  1417 => (x"fd",x"49",x"73",x"87"),
  1418 => (x"4b",x"26",x"87",x"f4"),
  1419 => (x"73",x"1e",x"4f",x"26"),
  1420 => (x"c2",x"4b",x"71",x"1e"),
  1421 => (x"d6",x"02",x"4a",x"a3"),
  1422 => (x"05",x"8a",x"c1",x"87"),
  1423 => (x"c2",x"87",x"e2",x"c0"),
  1424 => (x"02",x"bf",x"d8",x"f4"),
  1425 => (x"c1",x"48",x"87",x"db"),
  1426 => (x"dc",x"f4",x"c2",x"88"),
  1427 => (x"c2",x"87",x"d2",x"58"),
  1428 => (x"02",x"bf",x"dc",x"f4"),
  1429 => (x"f4",x"c2",x"87",x"cb"),
  1430 => (x"c1",x"48",x"bf",x"d8"),
  1431 => (x"dc",x"f4",x"c2",x"80"),
  1432 => (x"c2",x"1e",x"c7",x"58"),
  1433 => (x"1e",x"bf",x"d8",x"f4"),
  1434 => (x"1e",x"ec",x"ed",x"c1"),
  1435 => (x"97",x"c8",x"f3",x"c2"),
  1436 => (x"87",x"cc",x"49",x"bf"),
  1437 => (x"f2",x"c0",x"49",x"73"),
  1438 => (x"8e",x"f4",x"87",x"c6"),
  1439 => (x"4f",x"26",x"4b",x"26"),
  1440 => (x"5c",x"5b",x"5e",x"0e"),
  1441 => (x"cc",x"ff",x"0e",x"5d"),
  1442 => (x"a6",x"e8",x"c0",x"86"),
  1443 => (x"48",x"a6",x"cc",x"59"),
  1444 => (x"80",x"c4",x"78",x"c0"),
  1445 => (x"80",x"c4",x"78",x"c0"),
  1446 => (x"80",x"c4",x"78",x"c0"),
  1447 => (x"78",x"66",x"c8",x"c1"),
  1448 => (x"78",x"c1",x"80",x"c4"),
  1449 => (x"78",x"c1",x"80",x"c4"),
  1450 => (x"48",x"dc",x"f4",x"c2"),
  1451 => (x"df",x"ff",x"78",x"c1"),
  1452 => (x"c3",x"e0",x"87",x"e9"),
  1453 => (x"d7",x"df",x"ff",x"87"),
  1454 => (x"c0",x"4d",x"70",x"87"),
  1455 => (x"c1",x"02",x"ad",x"fb"),
  1456 => (x"e4",x"c0",x"87",x"f3"),
  1457 => (x"e8",x"c1",x"05",x"66"),
  1458 => (x"66",x"c4",x"c1",x"87"),
  1459 => (x"6a",x"82",x"c4",x"4a"),
  1460 => (x"d0",x"ca",x"c1",x"7e"),
  1461 => (x"20",x"49",x"6e",x"48"),
  1462 => (x"10",x"41",x"20",x"41"),
  1463 => (x"66",x"c4",x"c1",x"51"),
  1464 => (x"ca",x"d4",x"c1",x"48"),
  1465 => (x"c7",x"49",x"6a",x"78"),
  1466 => (x"c1",x"51",x"75",x"81"),
  1467 => (x"c8",x"49",x"66",x"c4"),
  1468 => (x"dc",x"51",x"c1",x"81"),
  1469 => (x"78",x"c2",x"48",x"a6"),
  1470 => (x"49",x"66",x"c4",x"c1"),
  1471 => (x"51",x"c0",x"81",x"c9"),
  1472 => (x"49",x"66",x"c4",x"c1"),
  1473 => (x"51",x"c0",x"81",x"ca"),
  1474 => (x"1e",x"d8",x"1e",x"c1"),
  1475 => (x"81",x"c8",x"49",x"6a"),
  1476 => (x"87",x"f8",x"de",x"ff"),
  1477 => (x"c8",x"c1",x"86",x"c8"),
  1478 => (x"a8",x"c0",x"48",x"66"),
  1479 => (x"d4",x"87",x"c7",x"01"),
  1480 => (x"78",x"c1",x"48",x"a6"),
  1481 => (x"c8",x"c1",x"87",x"cf"),
  1482 => (x"88",x"c1",x"48",x"66"),
  1483 => (x"c4",x"58",x"a6",x"dc"),
  1484 => (x"c3",x"de",x"ff",x"87"),
  1485 => (x"02",x"9d",x"75",x"87"),
  1486 => (x"d4",x"87",x"f1",x"cb"),
  1487 => (x"cc",x"c1",x"48",x"66"),
  1488 => (x"cb",x"03",x"a8",x"66"),
  1489 => (x"7e",x"c0",x"87",x"e6"),
  1490 => (x"87",x"c4",x"dd",x"ff"),
  1491 => (x"c1",x"48",x"4d",x"70"),
  1492 => (x"a6",x"c8",x"88",x"c6"),
  1493 => (x"02",x"98",x"70",x"58"),
  1494 => (x"48",x"87",x"d6",x"c1"),
  1495 => (x"a6",x"c8",x"88",x"c9"),
  1496 => (x"02",x"98",x"70",x"58"),
  1497 => (x"48",x"87",x"d7",x"c5"),
  1498 => (x"a6",x"c8",x"88",x"c1"),
  1499 => (x"02",x"98",x"70",x"58"),
  1500 => (x"48",x"87",x"f8",x"c2"),
  1501 => (x"a6",x"c8",x"88",x"c3"),
  1502 => (x"02",x"98",x"70",x"58"),
  1503 => (x"c1",x"48",x"87",x"cf"),
  1504 => (x"58",x"a6",x"c8",x"88"),
  1505 => (x"c4",x"02",x"98",x"70"),
  1506 => (x"fe",x"c9",x"87",x"f4"),
  1507 => (x"7e",x"f0",x"c0",x"87"),
  1508 => (x"87",x"fc",x"db",x"ff"),
  1509 => (x"ec",x"c0",x"4d",x"70"),
  1510 => (x"87",x"c2",x"02",x"ad"),
  1511 => (x"ec",x"c0",x"7e",x"75"),
  1512 => (x"87",x"cd",x"02",x"ad"),
  1513 => (x"87",x"e8",x"db",x"ff"),
  1514 => (x"ec",x"c0",x"4d",x"70"),
  1515 => (x"f3",x"ff",x"05",x"ad"),
  1516 => (x"66",x"e4",x"c0",x"87"),
  1517 => (x"87",x"ea",x"c1",x"05"),
  1518 => (x"02",x"ad",x"ec",x"c0"),
  1519 => (x"db",x"ff",x"87",x"c4"),
  1520 => (x"1e",x"c0",x"87",x"ce"),
  1521 => (x"66",x"dc",x"1e",x"ca"),
  1522 => (x"c1",x"93",x"cc",x"4b"),
  1523 => (x"c4",x"83",x"66",x"cc"),
  1524 => (x"49",x"6c",x"4c",x"a3"),
  1525 => (x"87",x"f4",x"db",x"ff"),
  1526 => (x"1e",x"de",x"1e",x"c1"),
  1527 => (x"db",x"ff",x"49",x"6c"),
  1528 => (x"86",x"d0",x"87",x"ea"),
  1529 => (x"7b",x"ca",x"d4",x"c1"),
  1530 => (x"dc",x"49",x"a3",x"c8"),
  1531 => (x"a3",x"c9",x"51",x"66"),
  1532 => (x"66",x"e0",x"c0",x"49"),
  1533 => (x"49",x"a3",x"ca",x"51"),
  1534 => (x"66",x"dc",x"51",x"6e"),
  1535 => (x"c0",x"80",x"c1",x"48"),
  1536 => (x"d4",x"58",x"a6",x"e0"),
  1537 => (x"66",x"d8",x"48",x"66"),
  1538 => (x"87",x"cb",x"04",x"a8"),
  1539 => (x"c1",x"48",x"66",x"d4"),
  1540 => (x"58",x"a6",x"d8",x"80"),
  1541 => (x"d8",x"87",x"fa",x"c7"),
  1542 => (x"88",x"c1",x"48",x"66"),
  1543 => (x"c7",x"58",x"a6",x"dc"),
  1544 => (x"da",x"ff",x"87",x"ef"),
  1545 => (x"4d",x"70",x"87",x"d2"),
  1546 => (x"ff",x"87",x"e6",x"c7"),
  1547 => (x"d0",x"87",x"c8",x"dc"),
  1548 => (x"66",x"d0",x"58",x"a6"),
  1549 => (x"87",x"c6",x"06",x"a8"),
  1550 => (x"cc",x"48",x"a6",x"d0"),
  1551 => (x"db",x"ff",x"78",x"66"),
  1552 => (x"ec",x"c0",x"87",x"f5"),
  1553 => (x"f5",x"c1",x"05",x"a8"),
  1554 => (x"66",x"e4",x"c0",x"87"),
  1555 => (x"87",x"e5",x"c1",x"05"),
  1556 => (x"cc",x"49",x"66",x"d4"),
  1557 => (x"66",x"c4",x"c1",x"91"),
  1558 => (x"4a",x"a1",x"c4",x"81"),
  1559 => (x"a1",x"c8",x"4c",x"6a"),
  1560 => (x"52",x"66",x"cc",x"4a"),
  1561 => (x"79",x"d0",x"d5",x"c1"),
  1562 => (x"87",x"e4",x"d8",x"ff"),
  1563 => (x"02",x"9d",x"4d",x"70"),
  1564 => (x"fb",x"c0",x"87",x"da"),
  1565 => (x"87",x"d4",x"02",x"ad"),
  1566 => (x"d8",x"ff",x"54",x"75"),
  1567 => (x"4d",x"70",x"87",x"d2"),
  1568 => (x"c7",x"c0",x"02",x"9d"),
  1569 => (x"ad",x"fb",x"c0",x"87"),
  1570 => (x"87",x"ec",x"ff",x"05"),
  1571 => (x"c2",x"54",x"e0",x"c0"),
  1572 => (x"97",x"c0",x"54",x"c1"),
  1573 => (x"48",x"66",x"d4",x"7c"),
  1574 => (x"04",x"a8",x"66",x"d8"),
  1575 => (x"d4",x"87",x"cb",x"c0"),
  1576 => (x"80",x"c1",x"48",x"66"),
  1577 => (x"c5",x"58",x"a6",x"d8"),
  1578 => (x"66",x"d8",x"87",x"e7"),
  1579 => (x"dc",x"88",x"c1",x"48"),
  1580 => (x"dc",x"c5",x"58",x"a6"),
  1581 => (x"ff",x"d7",x"ff",x"87"),
  1582 => (x"c5",x"4d",x"70",x"87"),
  1583 => (x"66",x"cc",x"87",x"d3"),
  1584 => (x"66",x"e4",x"c0",x"48"),
  1585 => (x"f4",x"c4",x"05",x"a8"),
  1586 => (x"a6",x"e8",x"c0",x"87"),
  1587 => (x"ff",x"78",x"c0",x"48"),
  1588 => (x"70",x"87",x"e4",x"d9"),
  1589 => (x"de",x"d9",x"ff",x"7e"),
  1590 => (x"a6",x"f0",x"c0",x"87"),
  1591 => (x"a8",x"ec",x"c0",x"58"),
  1592 => (x"87",x"c7",x"c0",x"05"),
  1593 => (x"78",x"6e",x"48",x"a6"),
  1594 => (x"ff",x"87",x"c4",x"c0"),
  1595 => (x"d4",x"87",x"e1",x"d6"),
  1596 => (x"91",x"cc",x"49",x"66"),
  1597 => (x"48",x"66",x"c4",x"c1"),
  1598 => (x"a6",x"c8",x"80",x"71"),
  1599 => (x"4a",x"66",x"c4",x"58"),
  1600 => (x"66",x"c4",x"82",x"c8"),
  1601 => (x"6e",x"81",x"ca",x"49"),
  1602 => (x"66",x"ec",x"c0",x"51"),
  1603 => (x"6e",x"81",x"c1",x"49"),
  1604 => (x"71",x"48",x"c1",x"89"),
  1605 => (x"c1",x"49",x"70",x"30"),
  1606 => (x"7a",x"97",x"71",x"89"),
  1607 => (x"bf",x"c4",x"f3",x"c2"),
  1608 => (x"97",x"29",x"6e",x"49"),
  1609 => (x"71",x"48",x"4a",x"6a"),
  1610 => (x"a6",x"f4",x"c0",x"98"),
  1611 => (x"48",x"66",x"c4",x"58"),
  1612 => (x"a6",x"cc",x"80",x"c4"),
  1613 => (x"bf",x"66",x"c8",x"58"),
  1614 => (x"66",x"e4",x"c0",x"4c"),
  1615 => (x"a8",x"66",x"cc",x"48"),
  1616 => (x"87",x"c5",x"c0",x"02"),
  1617 => (x"c2",x"c0",x"7e",x"c0"),
  1618 => (x"6e",x"7e",x"c1",x"87"),
  1619 => (x"1e",x"e0",x"c0",x"1e"),
  1620 => (x"d5",x"ff",x"49",x"74"),
  1621 => (x"86",x"c8",x"87",x"f6"),
  1622 => (x"b7",x"c0",x"4d",x"70"),
  1623 => (x"d4",x"c1",x"06",x"ad"),
  1624 => (x"c8",x"84",x"75",x"87"),
  1625 => (x"c0",x"49",x"bf",x"66"),
  1626 => (x"89",x"74",x"81",x"e0"),
  1627 => (x"dc",x"ca",x"c1",x"4b"),
  1628 => (x"de",x"fe",x"71",x"4a"),
  1629 => (x"84",x"c2",x"87",x"ed"),
  1630 => (x"e8",x"c0",x"7e",x"74"),
  1631 => (x"80",x"c1",x"48",x"66"),
  1632 => (x"58",x"a6",x"ec",x"c0"),
  1633 => (x"49",x"66",x"f0",x"c0"),
  1634 => (x"a9",x"70",x"81",x"c1"),
  1635 => (x"87",x"c5",x"c0",x"02"),
  1636 => (x"c2",x"c0",x"4c",x"c0"),
  1637 => (x"74",x"4c",x"c1",x"87"),
  1638 => (x"bf",x"66",x"cc",x"1e"),
  1639 => (x"81",x"e0",x"c0",x"49"),
  1640 => (x"71",x"89",x"66",x"c4"),
  1641 => (x"49",x"66",x"c8",x"1e"),
  1642 => (x"87",x"e0",x"d4",x"ff"),
  1643 => (x"b7",x"c0",x"86",x"c8"),
  1644 => (x"c5",x"ff",x"01",x"a8"),
  1645 => (x"66",x"e8",x"c0",x"87"),
  1646 => (x"87",x"d3",x"c0",x"02"),
  1647 => (x"c9",x"49",x"66",x"c4"),
  1648 => (x"66",x"e8",x"c0",x"81"),
  1649 => (x"48",x"66",x"c4",x"51"),
  1650 => (x"78",x"de",x"d6",x"c1"),
  1651 => (x"c4",x"87",x"ce",x"c0"),
  1652 => (x"81",x"c9",x"49",x"66"),
  1653 => (x"66",x"c4",x"51",x"c2"),
  1654 => (x"dc",x"d8",x"c1",x"48"),
  1655 => (x"48",x"66",x"d4",x"78"),
  1656 => (x"04",x"a8",x"66",x"d8"),
  1657 => (x"d4",x"87",x"cb",x"c0"),
  1658 => (x"80",x"c1",x"48",x"66"),
  1659 => (x"c0",x"58",x"a6",x"d8"),
  1660 => (x"66",x"d8",x"87",x"d1"),
  1661 => (x"dc",x"88",x"c1",x"48"),
  1662 => (x"c6",x"c0",x"58",x"a6"),
  1663 => (x"f7",x"d2",x"ff",x"87"),
  1664 => (x"cc",x"4d",x"70",x"87"),
  1665 => (x"78",x"c0",x"48",x"a6"),
  1666 => (x"ff",x"87",x"c6",x"c0"),
  1667 => (x"70",x"87",x"e9",x"d2"),
  1668 => (x"66",x"e0",x"c0",x"4d"),
  1669 => (x"c0",x"80",x"c1",x"48"),
  1670 => (x"75",x"58",x"a6",x"e4"),
  1671 => (x"cb",x"c0",x"02",x"9d"),
  1672 => (x"48",x"66",x"d4",x"87"),
  1673 => (x"a8",x"66",x"cc",x"c1"),
  1674 => (x"87",x"da",x"f4",x"04"),
  1675 => (x"c7",x"48",x"66",x"d4"),
  1676 => (x"e1",x"c0",x"03",x"a8"),
  1677 => (x"4c",x"66",x"d4",x"87"),
  1678 => (x"48",x"dc",x"f4",x"c2"),
  1679 => (x"49",x"74",x"78",x"c0"),
  1680 => (x"c4",x"c1",x"91",x"cc"),
  1681 => (x"a1",x"c4",x"81",x"66"),
  1682 => (x"c0",x"4a",x"6a",x"4a"),
  1683 => (x"84",x"c1",x"79",x"52"),
  1684 => (x"ff",x"04",x"ac",x"c7"),
  1685 => (x"e4",x"c0",x"87",x"e2"),
  1686 => (x"e2",x"c0",x"02",x"66"),
  1687 => (x"66",x"c4",x"c1",x"87"),
  1688 => (x"81",x"d4",x"c1",x"49"),
  1689 => (x"4a",x"66",x"c4",x"c1"),
  1690 => (x"c0",x"82",x"dc",x"c1"),
  1691 => (x"d0",x"d5",x"c1",x"52"),
  1692 => (x"66",x"c4",x"c1",x"79"),
  1693 => (x"81",x"d8",x"c1",x"49"),
  1694 => (x"79",x"e0",x"ca",x"c1"),
  1695 => (x"c1",x"87",x"d6",x"c0"),
  1696 => (x"c1",x"49",x"66",x"c4"),
  1697 => (x"c4",x"c1",x"81",x"d4"),
  1698 => (x"d8",x"c1",x"4a",x"66"),
  1699 => (x"e8",x"ca",x"c1",x"82"),
  1700 => (x"c7",x"d5",x"c1",x"7a"),
  1701 => (x"66",x"c4",x"c1",x"79"),
  1702 => (x"81",x"e0",x"c1",x"49"),
  1703 => (x"79",x"ee",x"d8",x"c1"),
  1704 => (x"87",x"cb",x"d0",x"ff"),
  1705 => (x"ff",x"48",x"66",x"d0"),
  1706 => (x"4d",x"26",x"8e",x"cc"),
  1707 => (x"4b",x"26",x"4c",x"26"),
  1708 => (x"c7",x"1e",x"4f",x"26"),
  1709 => (x"d8",x"f4",x"c2",x"1e"),
  1710 => (x"ed",x"c1",x"1e",x"bf"),
  1711 => (x"f3",x"c2",x"1e",x"ec"),
  1712 => (x"49",x"bf",x"97",x"c8"),
  1713 => (x"c1",x"87",x"f9",x"ee"),
  1714 => (x"c0",x"49",x"ec",x"ed"),
  1715 => (x"f4",x"87",x"ff",x"e1"),
  1716 => (x"1e",x"4f",x"26",x"8e"),
  1717 => (x"48",x"e0",x"ed",x"c1"),
  1718 => (x"ef",x"c1",x"50",x"c0"),
  1719 => (x"ff",x"49",x"bf",x"d8"),
  1720 => (x"c0",x"87",x"c3",x"d5"),
  1721 => (x"1e",x"4f",x"26",x"48"),
  1722 => (x"cd",x"c7",x"1e",x"73"),
  1723 => (x"e4",x"f4",x"c2",x"87"),
  1724 => (x"ff",x"50",x"c0",x"48"),
  1725 => (x"ff",x"c3",x"48",x"d4"),
  1726 => (x"f0",x"ca",x"c1",x"78"),
  1727 => (x"e6",x"d6",x"fe",x"49"),
  1728 => (x"db",x"e2",x"fe",x"87"),
  1729 => (x"02",x"98",x"70",x"87"),
  1730 => (x"eb",x"fe",x"87",x"cd"),
  1731 => (x"98",x"70",x"87",x"f9"),
  1732 => (x"c1",x"87",x"c4",x"02"),
  1733 => (x"c0",x"87",x"c2",x"4a"),
  1734 => (x"02",x"9a",x"72",x"4a"),
  1735 => (x"ca",x"c1",x"87",x"c8"),
  1736 => (x"d6",x"fe",x"49",x"fc"),
  1737 => (x"f4",x"c2",x"87",x"c1"),
  1738 => (x"78",x"c0",x"48",x"d8"),
  1739 => (x"48",x"c8",x"f3",x"c2"),
  1740 => (x"fd",x"49",x"50",x"c0"),
  1741 => (x"da",x"fe",x"87",x"fc"),
  1742 => (x"9b",x"4b",x"70",x"87"),
  1743 => (x"c1",x"87",x"cf",x"02"),
  1744 => (x"c7",x"5b",x"c8",x"ef"),
  1745 => (x"87",x"f8",x"de",x"49"),
  1746 => (x"e0",x"c0",x"49",x"c1"),
  1747 => (x"f2",x"c2",x"87",x"d3"),
  1748 => (x"f4",x"e1",x"c0",x"87"),
  1749 => (x"d0",x"f1",x"c0",x"87"),
  1750 => (x"87",x"f5",x"ff",x"87"),
  1751 => (x"4f",x"26",x"4b",x"26"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"01"),
  1755 => (x"00",x"00",x"11",x"fa"),
  1756 => (x"00",x"00",x"2d",x"30"),
  1757 => (x"94",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"11",x"fa"),
  1759 => (x"00",x"00",x"2d",x"4e"),
  1760 => (x"94",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"11",x"fa"),
  1762 => (x"00",x"00",x"2d",x"6c"),
  1763 => (x"94",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"11",x"fa"),
  1765 => (x"00",x"00",x"2d",x"8a"),
  1766 => (x"94",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"11",x"fa"),
  1768 => (x"00",x"00",x"2d",x"a8"),
  1769 => (x"94",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"11",x"fa"),
  1771 => (x"00",x"00",x"2d",x"c6"),
  1772 => (x"94",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"11",x"fa"),
  1774 => (x"00",x"00",x"2d",x"e4"),
  1775 => (x"94",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"15",x"50"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"94",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"12",x"f4"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"94",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"12",x"c0"),
  1783 => (x"db",x"86",x"fc",x"1e"),
  1784 => (x"fc",x"7e",x"70",x"87"),
  1785 => (x"1e",x"4f",x"26",x"8e"),
  1786 => (x"c0",x"48",x"f0",x"fe"),
  1787 => (x"79",x"09",x"cd",x"78"),
  1788 => (x"1e",x"4f",x"26",x"09"),
  1789 => (x"49",x"dc",x"ef",x"c1"),
  1790 => (x"4f",x"26",x"87",x"ed"),
  1791 => (x"bf",x"f0",x"fe",x"1e"),
  1792 => (x"1e",x"4f",x"26",x"48"),
  1793 => (x"c1",x"48",x"f0",x"fe"),
  1794 => (x"1e",x"4f",x"26",x"78"),
  1795 => (x"c0",x"48",x"f0",x"fe"),
  1796 => (x"1e",x"4f",x"26",x"78"),
  1797 => (x"52",x"c0",x"4a",x"71"),
  1798 => (x"0e",x"4f",x"26",x"51"),
  1799 => (x"5d",x"5c",x"5b",x"5e"),
  1800 => (x"71",x"86",x"f4",x"0e"),
  1801 => (x"7e",x"6d",x"97",x"4d"),
  1802 => (x"97",x"4c",x"a5",x"c1"),
  1803 => (x"a6",x"c8",x"48",x"6c"),
  1804 => (x"c4",x"48",x"6e",x"58"),
  1805 => (x"c5",x"05",x"a8",x"66"),
  1806 => (x"c0",x"48",x"ff",x"87"),
  1807 => (x"ca",x"ff",x"87",x"e6"),
  1808 => (x"49",x"a5",x"c2",x"87"),
  1809 => (x"71",x"4b",x"6c",x"97"),
  1810 => (x"6b",x"97",x"4b",x"a3"),
  1811 => (x"7e",x"6c",x"97",x"4b"),
  1812 => (x"80",x"c1",x"48",x"6e"),
  1813 => (x"c7",x"58",x"a6",x"c8"),
  1814 => (x"58",x"a6",x"cc",x"98"),
  1815 => (x"fe",x"7c",x"97",x"70"),
  1816 => (x"48",x"73",x"87",x"e1"),
  1817 => (x"4d",x"26",x"8e",x"f4"),
  1818 => (x"4b",x"26",x"4c",x"26"),
  1819 => (x"73",x"1e",x"4f",x"26"),
  1820 => (x"fe",x"86",x"f4",x"1e"),
  1821 => (x"bf",x"e0",x"87",x"d5"),
  1822 => (x"e0",x"c0",x"49",x"4b"),
  1823 => (x"c0",x"02",x"99",x"c0"),
  1824 => (x"4a",x"73",x"87",x"ea"),
  1825 => (x"c2",x"9a",x"ff",x"c3"),
  1826 => (x"bf",x"97",x"d8",x"f8"),
  1827 => (x"da",x"f8",x"c2",x"49"),
  1828 => (x"c2",x"51",x"72",x"81"),
  1829 => (x"bf",x"97",x"d8",x"f8"),
  1830 => (x"c1",x"48",x"6e",x"7e"),
  1831 => (x"58",x"a6",x"c8",x"80"),
  1832 => (x"a6",x"cc",x"98",x"c7"),
  1833 => (x"d8",x"f8",x"c2",x"58"),
  1834 => (x"50",x"66",x"c8",x"48"),
  1835 => (x"70",x"87",x"cd",x"fd"),
  1836 => (x"87",x"cf",x"fd",x"7e"),
  1837 => (x"4b",x"26",x"8e",x"f4"),
  1838 => (x"c2",x"1e",x"4f",x"26"),
  1839 => (x"fd",x"49",x"d8",x"f8"),
  1840 => (x"f1",x"c1",x"87",x"d1"),
  1841 => (x"de",x"fc",x"49",x"ee"),
  1842 => (x"87",x"e8",x"c4",x"87"),
  1843 => (x"5e",x"0e",x"4f",x"26"),
  1844 => (x"0e",x"5d",x"5c",x"5b"),
  1845 => (x"7e",x"71",x"86",x"fc"),
  1846 => (x"c2",x"4d",x"d4",x"ff"),
  1847 => (x"fc",x"49",x"d8",x"f8"),
  1848 => (x"4b",x"70",x"87",x"f9"),
  1849 => (x"04",x"ab",x"b7",x"c0"),
  1850 => (x"c3",x"87",x"f5",x"c2"),
  1851 => (x"c9",x"05",x"ab",x"f0"),
  1852 => (x"ec",x"f6",x"c1",x"87"),
  1853 => (x"c2",x"78",x"c1",x"48"),
  1854 => (x"e0",x"c3",x"87",x"d6"),
  1855 => (x"87",x"c9",x"05",x"ab"),
  1856 => (x"48",x"f0",x"f6",x"c1"),
  1857 => (x"c7",x"c2",x"78",x"c1"),
  1858 => (x"f0",x"f6",x"c1",x"87"),
  1859 => (x"87",x"c6",x"02",x"bf"),
  1860 => (x"4c",x"a3",x"c0",x"c2"),
  1861 => (x"4c",x"73",x"87",x"c2"),
  1862 => (x"bf",x"ec",x"f6",x"c1"),
  1863 => (x"87",x"e0",x"c0",x"02"),
  1864 => (x"b7",x"c4",x"49",x"74"),
  1865 => (x"f6",x"c1",x"91",x"29"),
  1866 => (x"4a",x"74",x"81",x"f4"),
  1867 => (x"92",x"c2",x"9a",x"cf"),
  1868 => (x"30",x"72",x"48",x"c1"),
  1869 => (x"ba",x"ff",x"4a",x"70"),
  1870 => (x"98",x"69",x"48",x"72"),
  1871 => (x"87",x"db",x"79",x"70"),
  1872 => (x"b7",x"c4",x"49",x"74"),
  1873 => (x"f6",x"c1",x"91",x"29"),
  1874 => (x"4a",x"74",x"81",x"f4"),
  1875 => (x"92",x"c2",x"9a",x"cf"),
  1876 => (x"30",x"72",x"48",x"c3"),
  1877 => (x"69",x"48",x"4a",x"70"),
  1878 => (x"6e",x"79",x"70",x"b0"),
  1879 => (x"87",x"e4",x"c0",x"05"),
  1880 => (x"c8",x"48",x"d0",x"ff"),
  1881 => (x"7d",x"c5",x"78",x"e1"),
  1882 => (x"bf",x"f0",x"f6",x"c1"),
  1883 => (x"c3",x"87",x"c3",x"02"),
  1884 => (x"f6",x"c1",x"7d",x"e0"),
  1885 => (x"c3",x"02",x"bf",x"ec"),
  1886 => (x"7d",x"f0",x"c3",x"87"),
  1887 => (x"d0",x"ff",x"7d",x"73"),
  1888 => (x"78",x"e0",x"c0",x"48"),
  1889 => (x"48",x"f0",x"f6",x"c1"),
  1890 => (x"f6",x"c1",x"78",x"c0"),
  1891 => (x"78",x"c0",x"48",x"ec"),
  1892 => (x"49",x"d8",x"f8",x"c2"),
  1893 => (x"70",x"87",x"c4",x"fa"),
  1894 => (x"ab",x"b7",x"c0",x"4b"),
  1895 => (x"87",x"cb",x"fd",x"03"),
  1896 => (x"8e",x"fc",x"48",x"c0"),
  1897 => (x"4c",x"26",x"4d",x"26"),
  1898 => (x"4f",x"26",x"4b",x"26"),
  1899 => (x"00",x"00",x"00",x"00"),
  1900 => (x"00",x"00",x"00",x"00"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"14",x"14",x"14",x"14"),
  1903 => (x"14",x"14",x"14",x"14"),
  1904 => (x"14",x"14",x"14",x"14"),
  1905 => (x"14",x"14",x"14",x"14"),
  1906 => (x"14",x"14",x"14",x"14"),
  1907 => (x"14",x"14",x"14",x"14"),
  1908 => (x"14",x"14",x"14",x"14"),
  1909 => (x"14",x"14",x"14",x"14"),
  1910 => (x"14",x"14",x"14",x"14"),
  1911 => (x"14",x"14",x"14",x"14"),
  1912 => (x"14",x"14",x"14",x"14"),
  1913 => (x"14",x"14",x"14",x"14"),
  1914 => (x"14",x"14",x"14",x"14"),
  1915 => (x"14",x"14",x"14",x"14"),
  1916 => (x"14",x"14",x"14",x"14"),
  1917 => (x"72",x"4a",x"c0",x"1e"),
  1918 => (x"c1",x"91",x"c4",x"49"),
  1919 => (x"c0",x"81",x"f4",x"f6"),
  1920 => (x"d0",x"82",x"c1",x"79"),
  1921 => (x"ee",x"04",x"aa",x"b7"),
  1922 => (x"0e",x"4f",x"26",x"87"),
  1923 => (x"5d",x"5c",x"5b",x"5e"),
  1924 => (x"f7",x"4d",x"71",x"0e"),
  1925 => (x"4a",x"75",x"87",x"f5"),
  1926 => (x"92",x"2a",x"b7",x"c4"),
  1927 => (x"82",x"f4",x"f6",x"c1"),
  1928 => (x"9c",x"cf",x"4c",x"75"),
  1929 => (x"49",x"6a",x"94",x"c2"),
  1930 => (x"c3",x"2b",x"74",x"4b"),
  1931 => (x"74",x"48",x"c2",x"9b"),
  1932 => (x"ff",x"4c",x"70",x"30"),
  1933 => (x"71",x"48",x"74",x"bc"),
  1934 => (x"f7",x"7a",x"70",x"98"),
  1935 => (x"48",x"73",x"87",x"c5"),
  1936 => (x"4c",x"26",x"4d",x"26"),
  1937 => (x"4f",x"26",x"4b",x"26"),
  1938 => (x"48",x"d0",x"ff",x"1e"),
  1939 => (x"71",x"78",x"e1",x"c8"),
  1940 => (x"08",x"d4",x"ff",x"48"),
  1941 => (x"1e",x"4f",x"26",x"78"),
  1942 => (x"c8",x"48",x"d0",x"ff"),
  1943 => (x"48",x"71",x"78",x"e1"),
  1944 => (x"78",x"08",x"d4",x"ff"),
  1945 => (x"ff",x"48",x"66",x"c4"),
  1946 => (x"26",x"78",x"08",x"d4"),
  1947 => (x"4a",x"71",x"1e",x"4f"),
  1948 => (x"1e",x"49",x"66",x"c4"),
  1949 => (x"de",x"ff",x"49",x"72"),
  1950 => (x"48",x"d0",x"ff",x"87"),
  1951 => (x"fc",x"78",x"e0",x"c0"),
  1952 => (x"1e",x"4f",x"26",x"8e"),
  1953 => (x"4a",x"71",x"1e",x"73"),
  1954 => (x"ab",x"b7",x"c2",x"4b"),
  1955 => (x"a3",x"87",x"c8",x"03"),
  1956 => (x"ff",x"c3",x"4a",x"49"),
  1957 => (x"ce",x"87",x"c7",x"9a"),
  1958 => (x"c3",x"4a",x"49",x"a3"),
  1959 => (x"66",x"c8",x"9a",x"ff"),
  1960 => (x"49",x"72",x"1e",x"49"),
  1961 => (x"fc",x"87",x"c6",x"ff"),
  1962 => (x"26",x"4b",x"26",x"8e"),
  1963 => (x"d0",x"ff",x"1e",x"4f"),
  1964 => (x"78",x"c9",x"c8",x"48"),
  1965 => (x"d4",x"ff",x"48",x"71"),
  1966 => (x"4f",x"26",x"78",x"08"),
  1967 => (x"49",x"4a",x"71",x"1e"),
  1968 => (x"d0",x"ff",x"87",x"eb"),
  1969 => (x"26",x"78",x"c8",x"48"),
  1970 => (x"1e",x"73",x"1e",x"4f"),
  1971 => (x"f8",x"c2",x"4b",x"71"),
  1972 => (x"c3",x"02",x"bf",x"f0"),
  1973 => (x"87",x"eb",x"c2",x"87"),
  1974 => (x"c8",x"48",x"d0",x"ff"),
  1975 => (x"48",x"73",x"78",x"c9"),
  1976 => (x"ff",x"b0",x"e0",x"c0"),
  1977 => (x"c2",x"78",x"08",x"d4"),
  1978 => (x"c0",x"48",x"e4",x"f8"),
  1979 => (x"02",x"66",x"c8",x"78"),
  1980 => (x"ff",x"c3",x"87",x"c5"),
  1981 => (x"c0",x"87",x"c2",x"49"),
  1982 => (x"ec",x"f8",x"c2",x"49"),
  1983 => (x"02",x"66",x"cc",x"59"),
  1984 => (x"d5",x"c5",x"87",x"c6"),
  1985 => (x"87",x"c4",x"4a",x"d5"),
  1986 => (x"4a",x"ff",x"ff",x"cf"),
  1987 => (x"5a",x"f0",x"f8",x"c2"),
  1988 => (x"48",x"f0",x"f8",x"c2"),
  1989 => (x"4b",x"26",x"78",x"c1"),
  1990 => (x"5e",x"0e",x"4f",x"26"),
  1991 => (x"0e",x"5d",x"5c",x"5b"),
  1992 => (x"f8",x"c2",x"4d",x"71"),
  1993 => (x"75",x"4b",x"bf",x"ec"),
  1994 => (x"87",x"cb",x"02",x"9d"),
  1995 => (x"c1",x"91",x"c8",x"49"),
  1996 => (x"71",x"4a",x"c0",x"fb"),
  1997 => (x"c1",x"87",x"c4",x"82"),
  1998 => (x"c0",x"4a",x"c0",x"ff"),
  1999 => (x"73",x"49",x"12",x"4c"),
  2000 => (x"e8",x"f8",x"c2",x"99"),
  2001 => (x"b8",x"71",x"48",x"bf"),
  2002 => (x"78",x"08",x"d4",x"ff"),
  2003 => (x"84",x"2b",x"b7",x"c1"),
  2004 => (x"04",x"ac",x"b7",x"c8"),
  2005 => (x"f8",x"c2",x"87",x"e7"),
  2006 => (x"c8",x"48",x"bf",x"e4"),
  2007 => (x"e8",x"f8",x"c2",x"80"),
  2008 => (x"26",x"4d",x"26",x"58"),
  2009 => (x"26",x"4b",x"26",x"4c"),
  2010 => (x"1e",x"73",x"1e",x"4f"),
  2011 => (x"4a",x"13",x"4b",x"71"),
  2012 => (x"87",x"cb",x"02",x"9a"),
  2013 => (x"e1",x"fe",x"49",x"72"),
  2014 => (x"9a",x"4a",x"13",x"87"),
  2015 => (x"26",x"87",x"f5",x"05"),
  2016 => (x"1e",x"4f",x"26",x"4b"),
  2017 => (x"bf",x"e4",x"f8",x"c2"),
  2018 => (x"e4",x"f8",x"c2",x"49"),
  2019 => (x"78",x"a1",x"c1",x"48"),
  2020 => (x"a9",x"b7",x"c0",x"c4"),
  2021 => (x"ff",x"87",x"db",x"03"),
  2022 => (x"f8",x"c2",x"48",x"d4"),
  2023 => (x"c2",x"78",x"bf",x"e8"),
  2024 => (x"49",x"bf",x"e4",x"f8"),
  2025 => (x"48",x"e4",x"f8",x"c2"),
  2026 => (x"c4",x"78",x"a1",x"c1"),
  2027 => (x"04",x"a9",x"b7",x"c0"),
  2028 => (x"d0",x"ff",x"87",x"e5"),
  2029 => (x"c2",x"78",x"c8",x"48"),
  2030 => (x"c0",x"48",x"f0",x"f8"),
  2031 => (x"00",x"4f",x"26",x"78"),
  2032 => (x"00",x"00",x"00",x"00"),
  2033 => (x"00",x"00",x"00",x"00"),
  2034 => (x"5f",x"00",x"00",x"00"),
  2035 => (x"00",x"00",x"00",x"5f"),
  2036 => (x"00",x"03",x"03",x"00"),
  2037 => (x"00",x"00",x"03",x"03"),
  2038 => (x"14",x"7f",x"7f",x"14"),
  2039 => (x"00",x"14",x"7f",x"7f"),
  2040 => (x"6b",x"2e",x"24",x"00"),
  2041 => (x"00",x"12",x"3a",x"6b"),
  2042 => (x"18",x"36",x"6a",x"4c"),
  2043 => (x"00",x"32",x"56",x"6c"),
  2044 => (x"59",x"4f",x"7e",x"30"),
  2045 => (x"40",x"68",x"3a",x"77"),
  2046 => (x"07",x"04",x"00",x"00"),
  2047 => (x"00",x"00",x"00",x"03"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

