
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"f9",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c4",x"f9",x"c2"),
    14 => (x"48",x"d0",x"e6",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d7",x"e7"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"49",x"72"),
    82 => (x"c2",x"7c",x"71",x"99"),
    83 => (x"05",x"bf",x"d0",x"e6"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"c3",x"29",x"d8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"d0",x"49",x"66",x"d0"),
    90 => (x"99",x"ff",x"c3",x"29"),
    91 => (x"66",x"d0",x"7c",x"71"),
    92 => (x"c3",x"29",x"c8",x"49"),
    93 => (x"7c",x"71",x"99",x"ff"),
    94 => (x"c3",x"49",x"66",x"d0"),
    95 => (x"7c",x"71",x"99",x"ff"),
    96 => (x"29",x"d0",x"49",x"72"),
    97 => (x"71",x"99",x"ff",x"c3"),
    98 => (x"c9",x"4b",x"6c",x"7c"),
    99 => (x"c3",x"4d",x"ff",x"f0"),
   100 => (x"d0",x"05",x"ab",x"ff"),
   101 => (x"7c",x"ff",x"c3",x"87"),
   102 => (x"8d",x"c1",x"4b",x"6c"),
   103 => (x"c3",x"87",x"c6",x"02"),
   104 => (x"f0",x"02",x"ab",x"ff"),
   105 => (x"fe",x"48",x"73",x"87"),
   106 => (x"c0",x"1e",x"87",x"c7"),
   107 => (x"48",x"d4",x"ff",x"49"),
   108 => (x"c1",x"78",x"ff",x"c3"),
   109 => (x"b7",x"c8",x"c3",x"81"),
   110 => (x"87",x"f1",x"04",x"a9"),
   111 => (x"73",x"1e",x"4f",x"26"),
   112 => (x"c4",x"87",x"e7",x"1e"),
   113 => (x"c0",x"4b",x"df",x"f8"),
   114 => (x"f0",x"ff",x"c0",x"1e"),
   115 => (x"fd",x"49",x"f7",x"c1"),
   116 => (x"86",x"c4",x"87",x"e7"),
   117 => (x"c0",x"05",x"a8",x"c1"),
   118 => (x"d4",x"ff",x"87",x"ea"),
   119 => (x"78",x"ff",x"c3",x"48"),
   120 => (x"c0",x"c0",x"c0",x"c1"),
   121 => (x"c0",x"1e",x"c0",x"c0"),
   122 => (x"e9",x"c1",x"f0",x"e1"),
   123 => (x"87",x"c9",x"fd",x"49"),
   124 => (x"98",x"70",x"86",x"c4"),
   125 => (x"ff",x"87",x"ca",x"05"),
   126 => (x"ff",x"c3",x"48",x"d4"),
   127 => (x"cb",x"48",x"c1",x"78"),
   128 => (x"87",x"e6",x"fe",x"87"),
   129 => (x"fe",x"05",x"8b",x"c1"),
   130 => (x"48",x"c0",x"87",x"fd"),
   131 => (x"1e",x"87",x"e6",x"fc"),
   132 => (x"d4",x"ff",x"1e",x"73"),
   133 => (x"78",x"ff",x"c3",x"48"),
   134 => (x"1e",x"c0",x"4b",x"d3"),
   135 => (x"c1",x"f0",x"ff",x"c0"),
   136 => (x"d4",x"fc",x"49",x"c1"),
   137 => (x"70",x"86",x"c4",x"87"),
   138 => (x"87",x"ca",x"05",x"98"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"48",x"c1",x"78",x"ff"),
   141 => (x"f1",x"fd",x"87",x"cb"),
   142 => (x"05",x"8b",x"c1",x"87"),
   143 => (x"c0",x"87",x"db",x"ff"),
   144 => (x"87",x"f1",x"fb",x"48"),
   145 => (x"5c",x"5b",x"5e",x"0e"),
   146 => (x"4c",x"d4",x"ff",x"0e"),
   147 => (x"c6",x"87",x"db",x"fd"),
   148 => (x"e1",x"c0",x"1e",x"ea"),
   149 => (x"49",x"c8",x"c1",x"f0"),
   150 => (x"c4",x"87",x"de",x"fb"),
   151 => (x"02",x"a8",x"c1",x"86"),
   152 => (x"ea",x"fe",x"87",x"c8"),
   153 => (x"c1",x"48",x"c0",x"87"),
   154 => (x"da",x"fa",x"87",x"e2"),
   155 => (x"cf",x"49",x"70",x"87"),
   156 => (x"c6",x"99",x"ff",x"ff"),
   157 => (x"c8",x"02",x"a9",x"ea"),
   158 => (x"87",x"d3",x"fe",x"87"),
   159 => (x"cb",x"c1",x"48",x"c0"),
   160 => (x"7c",x"ff",x"c3",x"87"),
   161 => (x"fc",x"4b",x"f1",x"c0"),
   162 => (x"98",x"70",x"87",x"f4"),
   163 => (x"87",x"eb",x"c0",x"02"),
   164 => (x"ff",x"c0",x"1e",x"c0"),
   165 => (x"49",x"fa",x"c1",x"f0"),
   166 => (x"c4",x"87",x"de",x"fa"),
   167 => (x"05",x"98",x"70",x"86"),
   168 => (x"ff",x"c3",x"87",x"d9"),
   169 => (x"c3",x"49",x"6c",x"7c"),
   170 => (x"7c",x"7c",x"7c",x"ff"),
   171 => (x"99",x"c0",x"c1",x"7c"),
   172 => (x"c1",x"87",x"c4",x"02"),
   173 => (x"c0",x"87",x"d5",x"48"),
   174 => (x"c2",x"87",x"d1",x"48"),
   175 => (x"87",x"c4",x"05",x"ab"),
   176 => (x"87",x"c8",x"48",x"c0"),
   177 => (x"fe",x"05",x"8b",x"c1"),
   178 => (x"48",x"c0",x"87",x"fd"),
   179 => (x"1e",x"87",x"e4",x"f9"),
   180 => (x"e6",x"c2",x"1e",x"73"),
   181 => (x"78",x"c1",x"48",x"d0"),
   182 => (x"d0",x"ff",x"4b",x"c7"),
   183 => (x"fb",x"78",x"c2",x"48"),
   184 => (x"d0",x"ff",x"87",x"c8"),
   185 => (x"c0",x"78",x"c3",x"48"),
   186 => (x"d0",x"e5",x"c0",x"1e"),
   187 => (x"f9",x"49",x"c0",x"c1"),
   188 => (x"86",x"c4",x"87",x"c7"),
   189 => (x"c1",x"05",x"a8",x"c1"),
   190 => (x"ab",x"c2",x"4b",x"87"),
   191 => (x"c0",x"87",x"c5",x"05"),
   192 => (x"87",x"f9",x"c0",x"48"),
   193 => (x"ff",x"05",x"8b",x"c1"),
   194 => (x"f7",x"fc",x"87",x"d0"),
   195 => (x"d4",x"e6",x"c2",x"87"),
   196 => (x"05",x"98",x"70",x"58"),
   197 => (x"1e",x"c1",x"87",x"cd"),
   198 => (x"c1",x"f0",x"ff",x"c0"),
   199 => (x"d8",x"f8",x"49",x"d0"),
   200 => (x"ff",x"86",x"c4",x"87"),
   201 => (x"ff",x"c3",x"48",x"d4"),
   202 => (x"87",x"de",x"c4",x"78"),
   203 => (x"58",x"d8",x"e6",x"c2"),
   204 => (x"c2",x"48",x"d0",x"ff"),
   205 => (x"48",x"d4",x"ff",x"78"),
   206 => (x"c1",x"78",x"ff",x"c3"),
   207 => (x"87",x"f5",x"f7",x"48"),
   208 => (x"5c",x"5b",x"5e",x"0e"),
   209 => (x"4a",x"71",x"0e",x"5d"),
   210 => (x"ff",x"4d",x"ff",x"c3"),
   211 => (x"7c",x"75",x"4c",x"d4"),
   212 => (x"c4",x"48",x"d0",x"ff"),
   213 => (x"7c",x"75",x"78",x"c3"),
   214 => (x"ff",x"c0",x"1e",x"72"),
   215 => (x"49",x"d8",x"c1",x"f0"),
   216 => (x"c4",x"87",x"d6",x"f7"),
   217 => (x"02",x"98",x"70",x"86"),
   218 => (x"48",x"c1",x"87",x"c5"),
   219 => (x"75",x"87",x"f0",x"c0"),
   220 => (x"7c",x"fe",x"c3",x"7c"),
   221 => (x"d4",x"1e",x"c0",x"c8"),
   222 => (x"fa",x"f4",x"49",x"66"),
   223 => (x"75",x"86",x"c4",x"87"),
   224 => (x"75",x"7c",x"75",x"7c"),
   225 => (x"e0",x"da",x"d8",x"7c"),
   226 => (x"6c",x"7c",x"75",x"4b"),
   227 => (x"c5",x"05",x"99",x"49"),
   228 => (x"05",x"8b",x"c1",x"87"),
   229 => (x"7c",x"75",x"87",x"f3"),
   230 => (x"c2",x"48",x"d0",x"ff"),
   231 => (x"f6",x"48",x"c0",x"78"),
   232 => (x"5e",x"0e",x"87",x"cf"),
   233 => (x"0e",x"5d",x"5c",x"5b"),
   234 => (x"4c",x"c0",x"4b",x"71"),
   235 => (x"df",x"cd",x"ee",x"c5"),
   236 => (x"48",x"d4",x"ff",x"4a"),
   237 => (x"68",x"78",x"ff",x"c3"),
   238 => (x"a9",x"fe",x"c3",x"49"),
   239 => (x"87",x"fd",x"c0",x"05"),
   240 => (x"9b",x"73",x"4d",x"70"),
   241 => (x"d0",x"87",x"cc",x"02"),
   242 => (x"49",x"73",x"1e",x"66"),
   243 => (x"c4",x"87",x"cf",x"f4"),
   244 => (x"ff",x"87",x"d6",x"86"),
   245 => (x"d1",x"c4",x"48",x"d0"),
   246 => (x"7d",x"ff",x"c3",x"78"),
   247 => (x"c1",x"48",x"66",x"d0"),
   248 => (x"58",x"a6",x"d4",x"88"),
   249 => (x"f0",x"05",x"98",x"70"),
   250 => (x"48",x"d4",x"ff",x"87"),
   251 => (x"78",x"78",x"ff",x"c3"),
   252 => (x"c5",x"05",x"9b",x"73"),
   253 => (x"48",x"d0",x"ff",x"87"),
   254 => (x"4a",x"c1",x"78",x"d0"),
   255 => (x"05",x"8a",x"c1",x"4c"),
   256 => (x"74",x"87",x"ee",x"fe"),
   257 => (x"87",x"e9",x"f4",x"48"),
   258 => (x"71",x"1e",x"73",x"1e"),
   259 => (x"ff",x"4b",x"c0",x"4a"),
   260 => (x"ff",x"c3",x"48",x"d4"),
   261 => (x"48",x"d0",x"ff",x"78"),
   262 => (x"ff",x"78",x"c3",x"c4"),
   263 => (x"ff",x"c3",x"48",x"d4"),
   264 => (x"c0",x"1e",x"72",x"78"),
   265 => (x"d1",x"c1",x"f0",x"ff"),
   266 => (x"87",x"cd",x"f4",x"49"),
   267 => (x"98",x"70",x"86",x"c4"),
   268 => (x"c8",x"87",x"d2",x"05"),
   269 => (x"66",x"cc",x"1e",x"c0"),
   270 => (x"87",x"e6",x"fd",x"49"),
   271 => (x"4b",x"70",x"86",x"c4"),
   272 => (x"c2",x"48",x"d0",x"ff"),
   273 => (x"f3",x"48",x"73",x"78"),
   274 => (x"5e",x"0e",x"87",x"eb"),
   275 => (x"0e",x"5d",x"5c",x"5b"),
   276 => (x"ff",x"c0",x"1e",x"c0"),
   277 => (x"49",x"c9",x"c1",x"f0"),
   278 => (x"d2",x"87",x"de",x"f3"),
   279 => (x"d8",x"e6",x"c2",x"1e"),
   280 => (x"87",x"fe",x"fc",x"49"),
   281 => (x"4c",x"c0",x"86",x"c8"),
   282 => (x"b7",x"d2",x"84",x"c1"),
   283 => (x"87",x"f8",x"04",x"ac"),
   284 => (x"97",x"d8",x"e6",x"c2"),
   285 => (x"c0",x"c3",x"49",x"bf"),
   286 => (x"a9",x"c0",x"c1",x"99"),
   287 => (x"87",x"e7",x"c0",x"05"),
   288 => (x"97",x"df",x"e6",x"c2"),
   289 => (x"31",x"d0",x"49",x"bf"),
   290 => (x"97",x"e0",x"e6",x"c2"),
   291 => (x"32",x"c8",x"4a",x"bf"),
   292 => (x"e6",x"c2",x"b1",x"72"),
   293 => (x"4a",x"bf",x"97",x"e1"),
   294 => (x"cf",x"4c",x"71",x"b1"),
   295 => (x"9c",x"ff",x"ff",x"ff"),
   296 => (x"34",x"ca",x"84",x"c1"),
   297 => (x"c2",x"87",x"e7",x"c1"),
   298 => (x"bf",x"97",x"e1",x"e6"),
   299 => (x"c6",x"31",x"c1",x"49"),
   300 => (x"e2",x"e6",x"c2",x"99"),
   301 => (x"c7",x"4a",x"bf",x"97"),
   302 => (x"b1",x"72",x"2a",x"b7"),
   303 => (x"97",x"dd",x"e6",x"c2"),
   304 => (x"cf",x"4d",x"4a",x"bf"),
   305 => (x"de",x"e6",x"c2",x"9d"),
   306 => (x"c3",x"4a",x"bf",x"97"),
   307 => (x"c2",x"32",x"ca",x"9a"),
   308 => (x"bf",x"97",x"df",x"e6"),
   309 => (x"73",x"33",x"c2",x"4b"),
   310 => (x"e0",x"e6",x"c2",x"b2"),
   311 => (x"c3",x"4b",x"bf",x"97"),
   312 => (x"b7",x"c6",x"9b",x"c0"),
   313 => (x"c2",x"b2",x"73",x"2b"),
   314 => (x"71",x"48",x"c1",x"81"),
   315 => (x"c1",x"49",x"70",x"30"),
   316 => (x"70",x"30",x"75",x"48"),
   317 => (x"c1",x"4c",x"72",x"4d"),
   318 => (x"c8",x"94",x"71",x"84"),
   319 => (x"06",x"ad",x"b7",x"c0"),
   320 => (x"34",x"c1",x"87",x"cc"),
   321 => (x"c0",x"c8",x"2d",x"b7"),
   322 => (x"ff",x"01",x"ad",x"b7"),
   323 => (x"48",x"74",x"87",x"f4"),
   324 => (x"0e",x"87",x"de",x"f0"),
   325 => (x"5d",x"5c",x"5b",x"5e"),
   326 => (x"c2",x"86",x"f8",x"0e"),
   327 => (x"c0",x"48",x"fe",x"ee"),
   328 => (x"f6",x"e6",x"c2",x"78"),
   329 => (x"fb",x"49",x"c0",x"1e"),
   330 => (x"86",x"c4",x"87",x"de"),
   331 => (x"c5",x"05",x"98",x"70"),
   332 => (x"c9",x"48",x"c0",x"87"),
   333 => (x"4d",x"c0",x"87",x"ce"),
   334 => (x"f2",x"c0",x"7e",x"c1"),
   335 => (x"c2",x"49",x"bf",x"ed"),
   336 => (x"71",x"4a",x"ec",x"e7"),
   337 => (x"e0",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"7e",x"c0",x"87",x"c2"),
   340 => (x"bf",x"e9",x"f2",x"c0"),
   341 => (x"c8",x"e8",x"c2",x"49"),
   342 => (x"4b",x"c8",x"71",x"4a"),
   343 => (x"70",x"87",x"ca",x"ec"),
   344 => (x"87",x"c2",x"05",x"98"),
   345 => (x"02",x"6e",x"7e",x"c0"),
   346 => (x"c2",x"87",x"fd",x"c0"),
   347 => (x"4d",x"bf",x"fc",x"ed"),
   348 => (x"9f",x"f4",x"ee",x"c2"),
   349 => (x"c5",x"48",x"7e",x"bf"),
   350 => (x"05",x"a8",x"ea",x"d6"),
   351 => (x"ed",x"c2",x"87",x"c7"),
   352 => (x"ce",x"4d",x"bf",x"fc"),
   353 => (x"ca",x"48",x"6e",x"87"),
   354 => (x"02",x"a8",x"d5",x"e9"),
   355 => (x"48",x"c0",x"87",x"c5"),
   356 => (x"c2",x"87",x"f1",x"c7"),
   357 => (x"75",x"1e",x"f6",x"e6"),
   358 => (x"87",x"ec",x"f9",x"49"),
   359 => (x"98",x"70",x"86",x"c4"),
   360 => (x"c0",x"87",x"c5",x"05"),
   361 => (x"87",x"dc",x"c7",x"48"),
   362 => (x"bf",x"e9",x"f2",x"c0"),
   363 => (x"c8",x"e8",x"c2",x"49"),
   364 => (x"4b",x"c8",x"71",x"4a"),
   365 => (x"70",x"87",x"f2",x"ea"),
   366 => (x"87",x"c8",x"05",x"98"),
   367 => (x"48",x"fe",x"ee",x"c2"),
   368 => (x"87",x"da",x"78",x"c1"),
   369 => (x"bf",x"ed",x"f2",x"c0"),
   370 => (x"ec",x"e7",x"c2",x"49"),
   371 => (x"4b",x"c8",x"71",x"4a"),
   372 => (x"70",x"87",x"d6",x"ea"),
   373 => (x"c5",x"c0",x"02",x"98"),
   374 => (x"c6",x"48",x"c0",x"87"),
   375 => (x"ee",x"c2",x"87",x"e6"),
   376 => (x"49",x"bf",x"97",x"f4"),
   377 => (x"05",x"a9",x"d5",x"c1"),
   378 => (x"c2",x"87",x"cd",x"c0"),
   379 => (x"bf",x"97",x"f5",x"ee"),
   380 => (x"a9",x"ea",x"c2",x"49"),
   381 => (x"87",x"c5",x"c0",x"02"),
   382 => (x"c7",x"c6",x"48",x"c0"),
   383 => (x"f6",x"e6",x"c2",x"87"),
   384 => (x"48",x"7e",x"bf",x"97"),
   385 => (x"02",x"a8",x"e9",x"c3"),
   386 => (x"6e",x"87",x"ce",x"c0"),
   387 => (x"a8",x"eb",x"c3",x"48"),
   388 => (x"87",x"c5",x"c0",x"02"),
   389 => (x"eb",x"c5",x"48",x"c0"),
   390 => (x"c1",x"e7",x"c2",x"87"),
   391 => (x"99",x"49",x"bf",x"97"),
   392 => (x"87",x"cc",x"c0",x"05"),
   393 => (x"97",x"c2",x"e7",x"c2"),
   394 => (x"a9",x"c2",x"49",x"bf"),
   395 => (x"87",x"c5",x"c0",x"02"),
   396 => (x"cf",x"c5",x"48",x"c0"),
   397 => (x"c3",x"e7",x"c2",x"87"),
   398 => (x"c2",x"48",x"bf",x"97"),
   399 => (x"70",x"58",x"fa",x"ee"),
   400 => (x"88",x"c1",x"48",x"4c"),
   401 => (x"58",x"fe",x"ee",x"c2"),
   402 => (x"97",x"c4",x"e7",x"c2"),
   403 => (x"81",x"75",x"49",x"bf"),
   404 => (x"97",x"c5",x"e7",x"c2"),
   405 => (x"32",x"c8",x"4a",x"bf"),
   406 => (x"c2",x"7e",x"a1",x"72"),
   407 => (x"6e",x"48",x"cb",x"f3"),
   408 => (x"c6",x"e7",x"c2",x"78"),
   409 => (x"c8",x"48",x"bf",x"97"),
   410 => (x"ee",x"c2",x"58",x"a6"),
   411 => (x"c2",x"02",x"bf",x"fe"),
   412 => (x"f2",x"c0",x"87",x"d4"),
   413 => (x"c2",x"49",x"bf",x"e9"),
   414 => (x"71",x"4a",x"c8",x"e8"),
   415 => (x"e8",x"e7",x"4b",x"c8"),
   416 => (x"02",x"98",x"70",x"87"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"f8",x"c3",x"48"),
   419 => (x"bf",x"f6",x"ee",x"c2"),
   420 => (x"df",x"f3",x"c2",x"4c"),
   421 => (x"db",x"e7",x"c2",x"5c"),
   422 => (x"c8",x"49",x"bf",x"97"),
   423 => (x"da",x"e7",x"c2",x"31"),
   424 => (x"a1",x"4a",x"bf",x"97"),
   425 => (x"dc",x"e7",x"c2",x"49"),
   426 => (x"d0",x"4a",x"bf",x"97"),
   427 => (x"49",x"a1",x"72",x"32"),
   428 => (x"97",x"dd",x"e7",x"c2"),
   429 => (x"32",x"d8",x"4a",x"bf"),
   430 => (x"c4",x"49",x"a1",x"72"),
   431 => (x"f3",x"c2",x"91",x"66"),
   432 => (x"c2",x"81",x"bf",x"cb"),
   433 => (x"c2",x"59",x"d3",x"f3"),
   434 => (x"bf",x"97",x"e3",x"e7"),
   435 => (x"c2",x"32",x"c8",x"4a"),
   436 => (x"bf",x"97",x"e2",x"e7"),
   437 => (x"c2",x"4a",x"a2",x"4b"),
   438 => (x"bf",x"97",x"e4",x"e7"),
   439 => (x"73",x"33",x"d0",x"4b"),
   440 => (x"e7",x"c2",x"4a",x"a2"),
   441 => (x"4b",x"bf",x"97",x"e5"),
   442 => (x"33",x"d8",x"9b",x"cf"),
   443 => (x"c2",x"4a",x"a2",x"73"),
   444 => (x"c2",x"5a",x"d7",x"f3"),
   445 => (x"4a",x"bf",x"d3",x"f3"),
   446 => (x"92",x"74",x"8a",x"c2"),
   447 => (x"48",x"d7",x"f3",x"c2"),
   448 => (x"c1",x"78",x"a1",x"72"),
   449 => (x"e7",x"c2",x"87",x"ca"),
   450 => (x"49",x"bf",x"97",x"c8"),
   451 => (x"e7",x"c2",x"31",x"c8"),
   452 => (x"4a",x"bf",x"97",x"c7"),
   453 => (x"ef",x"c2",x"49",x"a1"),
   454 => (x"ef",x"c2",x"59",x"c6"),
   455 => (x"c5",x"49",x"bf",x"c2"),
   456 => (x"81",x"ff",x"c7",x"31"),
   457 => (x"f3",x"c2",x"29",x"c9"),
   458 => (x"e7",x"c2",x"59",x"df"),
   459 => (x"4a",x"bf",x"97",x"cd"),
   460 => (x"e7",x"c2",x"32",x"c8"),
   461 => (x"4b",x"bf",x"97",x"cc"),
   462 => (x"66",x"c4",x"4a",x"a2"),
   463 => (x"c2",x"82",x"6e",x"92"),
   464 => (x"c2",x"5a",x"db",x"f3"),
   465 => (x"c0",x"48",x"d3",x"f3"),
   466 => (x"cf",x"f3",x"c2",x"78"),
   467 => (x"78",x"a1",x"72",x"48"),
   468 => (x"48",x"df",x"f3",x"c2"),
   469 => (x"bf",x"d3",x"f3",x"c2"),
   470 => (x"e3",x"f3",x"c2",x"78"),
   471 => (x"d7",x"f3",x"c2",x"48"),
   472 => (x"ee",x"c2",x"78",x"bf"),
   473 => (x"c0",x"02",x"bf",x"fe"),
   474 => (x"48",x"74",x"87",x"c9"),
   475 => (x"7e",x"70",x"30",x"c4"),
   476 => (x"c2",x"87",x"c9",x"c0"),
   477 => (x"48",x"bf",x"db",x"f3"),
   478 => (x"7e",x"70",x"30",x"c4"),
   479 => (x"48",x"c2",x"ef",x"c2"),
   480 => (x"48",x"c1",x"78",x"6e"),
   481 => (x"4d",x"26",x"8e",x"f8"),
   482 => (x"4b",x"26",x"4c",x"26"),
   483 => (x"5e",x"0e",x"4f",x"26"),
   484 => (x"0e",x"5d",x"5c",x"5b"),
   485 => (x"ee",x"c2",x"4a",x"71"),
   486 => (x"cb",x"02",x"bf",x"fe"),
   487 => (x"c7",x"4b",x"72",x"87"),
   488 => (x"c1",x"4c",x"72",x"2b"),
   489 => (x"87",x"c9",x"9c",x"ff"),
   490 => (x"2b",x"c8",x"4b",x"72"),
   491 => (x"ff",x"c3",x"4c",x"72"),
   492 => (x"cb",x"f3",x"c2",x"9c"),
   493 => (x"f2",x"c0",x"83",x"bf"),
   494 => (x"02",x"ab",x"bf",x"e5"),
   495 => (x"f2",x"c0",x"87",x"d9"),
   496 => (x"e6",x"c2",x"5b",x"e9"),
   497 => (x"49",x"73",x"1e",x"f6"),
   498 => (x"c4",x"87",x"fd",x"f0"),
   499 => (x"05",x"98",x"70",x"86"),
   500 => (x"48",x"c0",x"87",x"c5"),
   501 => (x"c2",x"87",x"e6",x"c0"),
   502 => (x"02",x"bf",x"fe",x"ee"),
   503 => (x"49",x"74",x"87",x"d2"),
   504 => (x"e6",x"c2",x"91",x"c4"),
   505 => (x"4d",x"69",x"81",x"f6"),
   506 => (x"ff",x"ff",x"ff",x"cf"),
   507 => (x"87",x"cb",x"9d",x"ff"),
   508 => (x"91",x"c2",x"49",x"74"),
   509 => (x"81",x"f6",x"e6",x"c2"),
   510 => (x"75",x"4d",x"69",x"9f"),
   511 => (x"87",x"c6",x"fe",x"48"),
   512 => (x"5c",x"5b",x"5e",x"0e"),
   513 => (x"86",x"f8",x"0e",x"5d"),
   514 => (x"05",x"9c",x"4c",x"71"),
   515 => (x"48",x"c0",x"87",x"c5"),
   516 => (x"c8",x"87",x"c2",x"c3"),
   517 => (x"48",x"6e",x"7e",x"a4"),
   518 => (x"66",x"d8",x"78",x"c0"),
   519 => (x"d8",x"87",x"c7",x"02"),
   520 => (x"05",x"bf",x"97",x"66"),
   521 => (x"48",x"c0",x"87",x"c5"),
   522 => (x"c0",x"87",x"ea",x"c2"),
   523 => (x"49",x"49",x"c1",x"1e"),
   524 => (x"c4",x"87",x"d7",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"c6",x"ef",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c8"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ed"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"d5",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"fe",x"ee"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ec"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"fa",x"ee",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fb",x"f9"),
   581 => (x"f6",x"ee",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"fa",x"ee",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d2",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"cf",x"f3",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"f6",x"ee",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"fa",x"ee",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"e9",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d5",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c7",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"cf",x"f3",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"f6",x"ee",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"fa",x"ee",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"e9"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"fe"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f8"),
   629 => (x"0e",x"5d",x"5c",x"5b"),
   630 => (x"d4",x"4b",x"71",x"1e"),
   631 => (x"9b",x"73",x"4d",x"66"),
   632 => (x"87",x"cc",x"c1",x"02"),
   633 => (x"69",x"49",x"a3",x"c8"),
   634 => (x"87",x"c4",x"c1",x"02"),
   635 => (x"c2",x"4c",x"a3",x"d0"),
   636 => (x"49",x"bf",x"fa",x"ee"),
   637 => (x"4a",x"6c",x"b9",x"ff"),
   638 => (x"66",x"d4",x"7e",x"99"),
   639 => (x"87",x"cd",x"06",x"a9"),
   640 => (x"cc",x"7c",x"7b",x"c0"),
   641 => (x"a3",x"c4",x"4a",x"a3"),
   642 => (x"ca",x"79",x"6a",x"49"),
   643 => (x"f8",x"49",x"72",x"87"),
   644 => (x"66",x"d4",x"99",x"c0"),
   645 => (x"75",x"8d",x"71",x"4d"),
   646 => (x"71",x"29",x"c9",x"49"),
   647 => (x"fa",x"49",x"73",x"1e"),
   648 => (x"e6",x"c2",x"87",x"f8"),
   649 => (x"49",x"73",x"1e",x"f6"),
   650 => (x"c8",x"87",x"c9",x"fc"),
   651 => (x"7c",x"66",x"d4",x"86"),
   652 => (x"87",x"d2",x"f5",x"26"),
   653 => (x"71",x"1e",x"73",x"1e"),
   654 => (x"c0",x"02",x"9b",x"4b"),
   655 => (x"f3",x"c2",x"87",x"e4"),
   656 => (x"4a",x"73",x"5b",x"e3"),
   657 => (x"ee",x"c2",x"8a",x"c2"),
   658 => (x"92",x"49",x"bf",x"f6"),
   659 => (x"bf",x"cf",x"f3",x"c2"),
   660 => (x"c2",x"80",x"72",x"48"),
   661 => (x"71",x"58",x"e7",x"f3"),
   662 => (x"c2",x"30",x"c4",x"48"),
   663 => (x"c0",x"58",x"c6",x"ef"),
   664 => (x"f3",x"c2",x"87",x"ed"),
   665 => (x"f3",x"c2",x"48",x"df"),
   666 => (x"c2",x"78",x"bf",x"d3"),
   667 => (x"c2",x"48",x"e3",x"f3"),
   668 => (x"78",x"bf",x"d7",x"f3"),
   669 => (x"bf",x"fe",x"ee",x"c2"),
   670 => (x"c2",x"87",x"c9",x"02"),
   671 => (x"49",x"bf",x"f6",x"ee"),
   672 => (x"87",x"c7",x"31",x"c4"),
   673 => (x"bf",x"db",x"f3",x"c2"),
   674 => (x"c2",x"31",x"c4",x"49"),
   675 => (x"f3",x"59",x"c6",x"ef"),
   676 => (x"5e",x"0e",x"87",x"f8"),
   677 => (x"71",x"0e",x"5c",x"5b"),
   678 => (x"72",x"4b",x"c0",x"4a"),
   679 => (x"e1",x"c0",x"02",x"9a"),
   680 => (x"49",x"a2",x"da",x"87"),
   681 => (x"c2",x"4b",x"69",x"9f"),
   682 => (x"02",x"bf",x"fe",x"ee"),
   683 => (x"a2",x"d4",x"87",x"cf"),
   684 => (x"49",x"69",x"9f",x"49"),
   685 => (x"ff",x"ff",x"c0",x"4c"),
   686 => (x"c2",x"34",x"d0",x"9c"),
   687 => (x"74",x"4c",x"c0",x"87"),
   688 => (x"49",x"73",x"b3",x"49"),
   689 => (x"f2",x"87",x"ed",x"fd"),
   690 => (x"5e",x"0e",x"87",x"fe"),
   691 => (x"0e",x"5d",x"5c",x"5b"),
   692 => (x"4a",x"71",x"86",x"f4"),
   693 => (x"9a",x"72",x"7e",x"c0"),
   694 => (x"c2",x"87",x"d8",x"02"),
   695 => (x"c0",x"48",x"f2",x"e6"),
   696 => (x"ea",x"e6",x"c2",x"78"),
   697 => (x"e3",x"f3",x"c2",x"48"),
   698 => (x"e6",x"c2",x"78",x"bf"),
   699 => (x"f3",x"c2",x"48",x"ee"),
   700 => (x"c2",x"78",x"bf",x"df"),
   701 => (x"c0",x"48",x"d3",x"ef"),
   702 => (x"c2",x"ef",x"c2",x"50"),
   703 => (x"e6",x"c2",x"49",x"bf"),
   704 => (x"71",x"4a",x"bf",x"f2"),
   705 => (x"c9",x"c4",x"03",x"aa"),
   706 => (x"cf",x"49",x"72",x"87"),
   707 => (x"e9",x"c0",x"05",x"99"),
   708 => (x"e5",x"f2",x"c0",x"87"),
   709 => (x"ea",x"e6",x"c2",x"48"),
   710 => (x"e6",x"c2",x"78",x"bf"),
   711 => (x"e6",x"c2",x"1e",x"f6"),
   712 => (x"c2",x"49",x"bf",x"ea"),
   713 => (x"c1",x"48",x"ea",x"e6"),
   714 => (x"e3",x"71",x"78",x"a1"),
   715 => (x"86",x"c4",x"87",x"da"),
   716 => (x"48",x"e1",x"f2",x"c0"),
   717 => (x"78",x"f6",x"e6",x"c2"),
   718 => (x"f2",x"c0",x"87",x"cc"),
   719 => (x"c0",x"48",x"bf",x"e1"),
   720 => (x"f2",x"c0",x"80",x"e0"),
   721 => (x"e6",x"c2",x"58",x"e5"),
   722 => (x"c1",x"48",x"bf",x"f2"),
   723 => (x"f6",x"e6",x"c2",x"80"),
   724 => (x"0c",x"a1",x"27",x"58"),
   725 => (x"97",x"bf",x"00",x"00"),
   726 => (x"02",x"9d",x"4d",x"bf"),
   727 => (x"c3",x"87",x"e3",x"c2"),
   728 => (x"c2",x"02",x"ad",x"e5"),
   729 => (x"f2",x"c0",x"87",x"dc"),
   730 => (x"cb",x"4b",x"bf",x"e1"),
   731 => (x"4c",x"11",x"49",x"a3"),
   732 => (x"c1",x"05",x"ac",x"cf"),
   733 => (x"49",x"75",x"87",x"d2"),
   734 => (x"89",x"c1",x"99",x"df"),
   735 => (x"ef",x"c2",x"91",x"cd"),
   736 => (x"a3",x"c1",x"81",x"c6"),
   737 => (x"c3",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"c5"),
   740 => (x"4a",x"a3",x"c7",x"51"),
   741 => (x"a3",x"c9",x"51",x"12"),
   742 => (x"ce",x"51",x"12",x"4a"),
   743 => (x"51",x"12",x"4a",x"a3"),
   744 => (x"12",x"4a",x"a3",x"d0"),
   745 => (x"4a",x"a3",x"d2",x"51"),
   746 => (x"a3",x"d4",x"51",x"12"),
   747 => (x"d6",x"51",x"12",x"4a"),
   748 => (x"51",x"12",x"4a",x"a3"),
   749 => (x"12",x"4a",x"a3",x"d8"),
   750 => (x"4a",x"a3",x"dc",x"51"),
   751 => (x"a3",x"de",x"51",x"12"),
   752 => (x"c1",x"51",x"12",x"4a"),
   753 => (x"87",x"fa",x"c0",x"7e"),
   754 => (x"99",x"c8",x"49",x"74"),
   755 => (x"87",x"eb",x"c0",x"05"),
   756 => (x"99",x"d0",x"49",x"74"),
   757 => (x"dc",x"87",x"d1",x"05"),
   758 => (x"cb",x"c0",x"02",x"66"),
   759 => (x"dc",x"49",x"73",x"87"),
   760 => (x"98",x"70",x"0f",x"66"),
   761 => (x"87",x"d3",x"c0",x"02"),
   762 => (x"c6",x"c0",x"05",x"6e"),
   763 => (x"c6",x"ef",x"c2",x"87"),
   764 => (x"c0",x"50",x"c0",x"48"),
   765 => (x"48",x"bf",x"e1",x"f2"),
   766 => (x"c2",x"87",x"e1",x"c2"),
   767 => (x"c0",x"48",x"d3",x"ef"),
   768 => (x"ef",x"c2",x"7e",x"50"),
   769 => (x"c2",x"49",x"bf",x"c2"),
   770 => (x"4a",x"bf",x"f2",x"e6"),
   771 => (x"fb",x"04",x"aa",x"71"),
   772 => (x"f3",x"c2",x"87",x"f7"),
   773 => (x"c0",x"05",x"bf",x"e3"),
   774 => (x"ee",x"c2",x"87",x"c8"),
   775 => (x"c1",x"02",x"bf",x"fe"),
   776 => (x"e6",x"c2",x"87",x"f8"),
   777 => (x"ed",x"49",x"bf",x"ee"),
   778 => (x"49",x"70",x"87",x"e4"),
   779 => (x"59",x"f2",x"e6",x"c2"),
   780 => (x"c2",x"48",x"a6",x"c4"),
   781 => (x"78",x"bf",x"ee",x"e6"),
   782 => (x"bf",x"fe",x"ee",x"c2"),
   783 => (x"87",x"d8",x"c0",x"02"),
   784 => (x"cf",x"49",x"66",x"c4"),
   785 => (x"f8",x"ff",x"ff",x"ff"),
   786 => (x"c0",x"02",x"a9",x"99"),
   787 => (x"4c",x"c0",x"87",x"c5"),
   788 => (x"c1",x"87",x"e1",x"c0"),
   789 => (x"87",x"dc",x"c0",x"4c"),
   790 => (x"cf",x"49",x"66",x"c4"),
   791 => (x"a9",x"99",x"f8",x"ff"),
   792 => (x"87",x"c8",x"c0",x"02"),
   793 => (x"c0",x"48",x"a6",x"c8"),
   794 => (x"87",x"c5",x"c0",x"78"),
   795 => (x"c1",x"48",x"a6",x"c8"),
   796 => (x"4c",x"66",x"c8",x"78"),
   797 => (x"c0",x"05",x"9c",x"74"),
   798 => (x"66",x"c4",x"87",x"e0"),
   799 => (x"c2",x"89",x"c2",x"49"),
   800 => (x"4a",x"bf",x"f6",x"ee"),
   801 => (x"cf",x"f3",x"c2",x"91"),
   802 => (x"e6",x"c2",x"4a",x"bf"),
   803 => (x"a1",x"72",x"48",x"ea"),
   804 => (x"f2",x"e6",x"c2",x"78"),
   805 => (x"f9",x"78",x"c0",x"48"),
   806 => (x"48",x"c0",x"87",x"df"),
   807 => (x"e5",x"eb",x"8e",x"f4"),
   808 => (x"00",x"00",x"00",x"87"),
   809 => (x"ff",x"ff",x"ff",x"00"),
   810 => (x"00",x"0c",x"b1",x"ff"),
   811 => (x"00",x"0c",x"ba",x"00"),
   812 => (x"54",x"41",x"46",x"00"),
   813 => (x"20",x"20",x"32",x"33"),
   814 => (x"41",x"46",x"00",x"20"),
   815 => (x"20",x"36",x"31",x"54"),
   816 => (x"1e",x"00",x"20",x"20"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"48",x"68",x"78",x"ff"),
   819 => (x"ff",x"1e",x"4f",x"26"),
   820 => (x"ff",x"c3",x"48",x"d4"),
   821 => (x"48",x"d0",x"ff",x"78"),
   822 => (x"ff",x"78",x"e1",x"c0"),
   823 => (x"78",x"d4",x"48",x"d4"),
   824 => (x"48",x"e7",x"f3",x"c2"),
   825 => (x"50",x"bf",x"d4",x"ff"),
   826 => (x"ff",x"1e",x"4f",x"26"),
   827 => (x"e0",x"c0",x"48",x"d0"),
   828 => (x"1e",x"4f",x"26",x"78"),
   829 => (x"70",x"87",x"cc",x"ff"),
   830 => (x"c6",x"02",x"99",x"49"),
   831 => (x"a9",x"fb",x"c0",x"87"),
   832 => (x"71",x"87",x"f1",x"05"),
   833 => (x"0e",x"4f",x"26",x"48"),
   834 => (x"0e",x"5c",x"5b",x"5e"),
   835 => (x"4c",x"c0",x"4b",x"71"),
   836 => (x"70",x"87",x"f0",x"fe"),
   837 => (x"c0",x"02",x"99",x"49"),
   838 => (x"ec",x"c0",x"87",x"f9"),
   839 => (x"f2",x"c0",x"02",x"a9"),
   840 => (x"a9",x"fb",x"c0",x"87"),
   841 => (x"87",x"eb",x"c0",x"02"),
   842 => (x"ac",x"b7",x"66",x"cc"),
   843 => (x"d0",x"87",x"c7",x"03"),
   844 => (x"87",x"c2",x"02",x"66"),
   845 => (x"99",x"71",x"53",x"71"),
   846 => (x"c1",x"87",x"c2",x"02"),
   847 => (x"87",x"c3",x"fe",x"84"),
   848 => (x"02",x"99",x"49",x"70"),
   849 => (x"ec",x"c0",x"87",x"cd"),
   850 => (x"87",x"c7",x"02",x"a9"),
   851 => (x"05",x"a9",x"fb",x"c0"),
   852 => (x"d0",x"87",x"d5",x"ff"),
   853 => (x"87",x"c3",x"02",x"66"),
   854 => (x"c0",x"7b",x"97",x"c0"),
   855 => (x"c4",x"05",x"a9",x"ec"),
   856 => (x"c5",x"4a",x"74",x"87"),
   857 => (x"c0",x"4a",x"74",x"87"),
   858 => (x"48",x"72",x"8a",x"0a"),
   859 => (x"4d",x"26",x"87",x"c2"),
   860 => (x"4b",x"26",x"4c",x"26"),
   861 => (x"fd",x"1e",x"4f",x"26"),
   862 => (x"49",x"70",x"87",x"c9"),
   863 => (x"aa",x"f0",x"c0",x"4a"),
   864 => (x"c0",x"87",x"c9",x"04"),
   865 => (x"c3",x"01",x"aa",x"f9"),
   866 => (x"8a",x"f0",x"c0",x"87"),
   867 => (x"04",x"aa",x"c1",x"c1"),
   868 => (x"da",x"c1",x"87",x"c9"),
   869 => (x"87",x"c3",x"01",x"aa"),
   870 => (x"72",x"8a",x"f7",x"c0"),
   871 => (x"0e",x"4f",x"26",x"48"),
   872 => (x"0e",x"5c",x"5b",x"5e"),
   873 => (x"d4",x"ff",x"4a",x"71"),
   874 => (x"c0",x"49",x"72",x"4b"),
   875 => (x"4c",x"70",x"87",x"e7"),
   876 => (x"87",x"c2",x"02",x"9c"),
   877 => (x"d0",x"ff",x"8c",x"c1"),
   878 => (x"c1",x"78",x"c5",x"48"),
   879 => (x"49",x"74",x"7b",x"d5"),
   880 => (x"e8",x"c1",x"31",x"c6"),
   881 => (x"4a",x"bf",x"97",x"f8"),
   882 => (x"70",x"b0",x"71",x"48"),
   883 => (x"48",x"d0",x"ff",x"7b"),
   884 => (x"db",x"fe",x"78",x"c4"),
   885 => (x"5b",x"5e",x"0e",x"87"),
   886 => (x"f8",x"0e",x"5d",x"5c"),
   887 => (x"c0",x"4b",x"71",x"86"),
   888 => (x"fc",x"fa",x"c0",x"7e"),
   889 => (x"df",x"49",x"bf",x"97"),
   890 => (x"ee",x"c0",x"05",x"a9"),
   891 => (x"49",x"a3",x"c8",x"87"),
   892 => (x"c1",x"49",x"69",x"97"),
   893 => (x"dd",x"05",x"a9",x"c3"),
   894 => (x"49",x"a3",x"c9",x"87"),
   895 => (x"c1",x"49",x"69",x"97"),
   896 => (x"d1",x"05",x"a9",x"c6"),
   897 => (x"49",x"a3",x"ca",x"87"),
   898 => (x"c1",x"49",x"69",x"97"),
   899 => (x"c5",x"05",x"a9",x"c7"),
   900 => (x"c2",x"48",x"c1",x"87"),
   901 => (x"48",x"c0",x"87",x"e1"),
   902 => (x"fa",x"87",x"dc",x"c2"),
   903 => (x"4c",x"c0",x"87",x"f0"),
   904 => (x"97",x"fc",x"fa",x"c0"),
   905 => (x"a9",x"c0",x"49",x"bf"),
   906 => (x"fb",x"87",x"cf",x"04"),
   907 => (x"84",x"c1",x"87",x"c5"),
   908 => (x"97",x"fc",x"fa",x"c0"),
   909 => (x"06",x"ac",x"49",x"bf"),
   910 => (x"fa",x"c0",x"87",x"f1"),
   911 => (x"02",x"bf",x"97",x"fc"),
   912 => (x"fe",x"f9",x"87",x"cf"),
   913 => (x"99",x"49",x"70",x"87"),
   914 => (x"c0",x"87",x"c6",x"02"),
   915 => (x"f1",x"05",x"a9",x"ec"),
   916 => (x"f9",x"4c",x"c0",x"87"),
   917 => (x"4d",x"70",x"87",x"ed"),
   918 => (x"c8",x"87",x"e8",x"f9"),
   919 => (x"e2",x"f9",x"58",x"a6"),
   920 => (x"c1",x"4a",x"70",x"87"),
   921 => (x"49",x"a3",x"c8",x"84"),
   922 => (x"ad",x"49",x"69",x"97"),
   923 => (x"c0",x"87",x"c7",x"02"),
   924 => (x"c0",x"05",x"ad",x"ff"),
   925 => (x"a3",x"c9",x"87",x"e7"),
   926 => (x"49",x"69",x"97",x"49"),
   927 => (x"02",x"a9",x"66",x"c4"),
   928 => (x"c0",x"48",x"87",x"c7"),
   929 => (x"d4",x"05",x"a8",x"ff"),
   930 => (x"49",x"a3",x"ca",x"87"),
   931 => (x"aa",x"49",x"69",x"97"),
   932 => (x"c0",x"87",x"c6",x"02"),
   933 => (x"c4",x"05",x"aa",x"ff"),
   934 => (x"d0",x"7e",x"c1",x"87"),
   935 => (x"ad",x"ec",x"c0",x"87"),
   936 => (x"c0",x"87",x"c6",x"02"),
   937 => (x"c4",x"05",x"ad",x"fb"),
   938 => (x"c1",x"4c",x"c0",x"87"),
   939 => (x"fe",x"02",x"6e",x"7e"),
   940 => (x"f5",x"f8",x"87",x"e1"),
   941 => (x"f8",x"48",x"74",x"87"),
   942 => (x"87",x"f2",x"fa",x"8e"),
   943 => (x"5b",x"5e",x"0e",x"00"),
   944 => (x"f8",x"0e",x"5d",x"5c"),
   945 => (x"ff",x"4d",x"71",x"86"),
   946 => (x"1e",x"75",x"4b",x"d4"),
   947 => (x"49",x"ec",x"f3",x"c2"),
   948 => (x"c4",x"87",x"ed",x"e4"),
   949 => (x"02",x"98",x"70",x"86"),
   950 => (x"c4",x"87",x"cc",x"c4"),
   951 => (x"e8",x"c1",x"48",x"a6"),
   952 => (x"75",x"78",x"bf",x"fa"),
   953 => (x"87",x"f7",x"fa",x"49"),
   954 => (x"c5",x"48",x"d0",x"ff"),
   955 => (x"7b",x"d6",x"c1",x"78"),
   956 => (x"a2",x"75",x"4a",x"c0"),
   957 => (x"c1",x"7b",x"11",x"49"),
   958 => (x"aa",x"b7",x"cb",x"82"),
   959 => (x"cc",x"87",x"f3",x"04"),
   960 => (x"7b",x"ff",x"c3",x"4a"),
   961 => (x"e0",x"c0",x"82",x"c1"),
   962 => (x"f4",x"04",x"aa",x"b7"),
   963 => (x"48",x"d0",x"ff",x"87"),
   964 => (x"ff",x"c3",x"78",x"c4"),
   965 => (x"c1",x"78",x"c5",x"7b"),
   966 => (x"7b",x"c1",x"7b",x"d3"),
   967 => (x"48",x"66",x"78",x"c4"),
   968 => (x"06",x"a8",x"b7",x"c0"),
   969 => (x"c2",x"87",x"f0",x"c2"),
   970 => (x"4c",x"bf",x"f4",x"f3"),
   971 => (x"74",x"48",x"66",x"c4"),
   972 => (x"58",x"a6",x"c8",x"88"),
   973 => (x"c1",x"02",x"9c",x"74"),
   974 => (x"e6",x"c2",x"87",x"f9"),
   975 => (x"c0",x"c8",x"7e",x"f6"),
   976 => (x"b7",x"c0",x"8c",x"4d"),
   977 => (x"87",x"c6",x"03",x"ac"),
   978 => (x"4d",x"a4",x"c0",x"c8"),
   979 => (x"f3",x"c2",x"4c",x"c0"),
   980 => (x"49",x"bf",x"97",x"e7"),
   981 => (x"d1",x"02",x"99",x"d0"),
   982 => (x"c2",x"1e",x"c0",x"87"),
   983 => (x"e7",x"49",x"ec",x"f3"),
   984 => (x"86",x"c4",x"87",x"d2"),
   985 => (x"c0",x"4a",x"49",x"70"),
   986 => (x"e6",x"c2",x"87",x"ee"),
   987 => (x"f3",x"c2",x"1e",x"f6"),
   988 => (x"ff",x"e6",x"49",x"ec"),
   989 => (x"70",x"86",x"c4",x"87"),
   990 => (x"d0",x"ff",x"4a",x"49"),
   991 => (x"78",x"c5",x"c8",x"48"),
   992 => (x"6e",x"7b",x"d4",x"c1"),
   993 => (x"6e",x"7b",x"bf",x"97"),
   994 => (x"70",x"80",x"c1",x"48"),
   995 => (x"05",x"8d",x"c1",x"7e"),
   996 => (x"ff",x"87",x"f0",x"ff"),
   997 => (x"78",x"c4",x"48",x"d0"),
   998 => (x"c5",x"05",x"9a",x"72"),
   999 => (x"c1",x"48",x"c0",x"87"),
  1000 => (x"1e",x"c1",x"87",x"c7"),
  1001 => (x"49",x"ec",x"f3",x"c2"),
  1002 => (x"c4",x"87",x"ef",x"e4"),
  1003 => (x"05",x"9c",x"74",x"86"),
  1004 => (x"c4",x"87",x"c7",x"fe"),
  1005 => (x"b7",x"c0",x"48",x"66"),
  1006 => (x"87",x"d1",x"06",x"a8"),
  1007 => (x"48",x"ec",x"f3",x"c2"),
  1008 => (x"80",x"d0",x"78",x"c0"),
  1009 => (x"80",x"f4",x"78",x"c0"),
  1010 => (x"bf",x"f8",x"f3",x"c2"),
  1011 => (x"48",x"66",x"c4",x"78"),
  1012 => (x"01",x"a8",x"b7",x"c0"),
  1013 => (x"ff",x"87",x"d0",x"fd"),
  1014 => (x"78",x"c5",x"48",x"d0"),
  1015 => (x"c0",x"7b",x"d3",x"c1"),
  1016 => (x"c1",x"78",x"c4",x"7b"),
  1017 => (x"c0",x"87",x"c2",x"48"),
  1018 => (x"26",x"8e",x"f8",x"48"),
  1019 => (x"26",x"4c",x"26",x"4d"),
  1020 => (x"0e",x"4f",x"26",x"4b"),
  1021 => (x"5d",x"5c",x"5b",x"5e"),
  1022 => (x"4b",x"71",x"1e",x"0e"),
  1023 => (x"ab",x"4d",x"4c",x"c0"),
  1024 => (x"87",x"e8",x"c0",x"04"),
  1025 => (x"1e",x"d5",x"f7",x"c0"),
  1026 => (x"c4",x"02",x"9d",x"75"),
  1027 => (x"c2",x"4a",x"c0",x"87"),
  1028 => (x"72",x"4a",x"c1",x"87"),
  1029 => (x"87",x"f2",x"ea",x"49"),
  1030 => (x"7e",x"70",x"86",x"c4"),
  1031 => (x"05",x"6e",x"84",x"c1"),
  1032 => (x"4c",x"73",x"87",x"c2"),
  1033 => (x"ac",x"73",x"85",x"c1"),
  1034 => (x"87",x"d8",x"ff",x"06"),
  1035 => (x"fe",x"26",x"48",x"6e"),
  1036 => (x"5e",x"0e",x"87",x"f9"),
  1037 => (x"71",x"0e",x"5c",x"5b"),
  1038 => (x"02",x"66",x"cc",x"4b"),
  1039 => (x"4c",x"87",x"e8",x"c0"),
  1040 => (x"02",x"8c",x"f0",x"c0"),
  1041 => (x"74",x"87",x"e8",x"c0"),
  1042 => (x"02",x"8a",x"c1",x"4a"),
  1043 => (x"8a",x"87",x"e0",x"c0"),
  1044 => (x"8a",x"87",x"dc",x"02"),
  1045 => (x"c0",x"87",x"d8",x"02"),
  1046 => (x"c0",x"02",x"8a",x"e0"),
  1047 => (x"8a",x"c1",x"87",x"e5"),
  1048 => (x"87",x"e7",x"c0",x"02"),
  1049 => (x"73",x"87",x"ea",x"c0"),
  1050 => (x"87",x"d1",x"f9",x"49"),
  1051 => (x"74",x"87",x"e2",x"c0"),
  1052 => (x"c1",x"49",x"c0",x"1e"),
  1053 => (x"74",x"87",x"f0",x"df"),
  1054 => (x"c1",x"49",x"73",x"1e"),
  1055 => (x"c8",x"87",x"e8",x"df"),
  1056 => (x"73",x"87",x"ce",x"86"),
  1057 => (x"d3",x"e2",x"c1",x"49"),
  1058 => (x"73",x"87",x"c6",x"87"),
  1059 => (x"c3",x"e3",x"c1",x"49"),
  1060 => (x"87",x"d9",x"fd",x"87"),
  1061 => (x"5c",x"5b",x"5e",x"0e"),
  1062 => (x"71",x"1e",x"0e",x"5d"),
  1063 => (x"91",x"de",x"49",x"4c"),
  1064 => (x"4d",x"d4",x"f4",x"c2"),
  1065 => (x"6d",x"97",x"85",x"71"),
  1066 => (x"87",x"de",x"c1",x"02"),
  1067 => (x"bf",x"c0",x"f4",x"c2"),
  1068 => (x"72",x"82",x"74",x"4a"),
  1069 => (x"87",x"fb",x"fc",x"49"),
  1070 => (x"98",x"48",x"7e",x"70"),
  1071 => (x"87",x"f2",x"c0",x"02"),
  1072 => (x"4b",x"c8",x"f4",x"c2"),
  1073 => (x"49",x"cb",x"4a",x"70"),
  1074 => (x"87",x"db",x"ff",x"fe"),
  1075 => (x"93",x"cb",x"4b",x"74"),
  1076 => (x"83",x"ef",x"e9",x"c1"),
  1077 => (x"c4",x"c1",x"83",x"c4"),
  1078 => (x"49",x"74",x"7b",x"ce"),
  1079 => (x"87",x"f0",x"c5",x"c1"),
  1080 => (x"e8",x"c1",x"7b",x"75"),
  1081 => (x"49",x"bf",x"97",x"f9"),
  1082 => (x"c8",x"f4",x"c2",x"1e"),
  1083 => (x"87",x"c2",x"fd",x"49"),
  1084 => (x"49",x"74",x"86",x"c4"),
  1085 => (x"87",x"d8",x"c5",x"c1"),
  1086 => (x"c6",x"c1",x"49",x"c0"),
  1087 => (x"f3",x"c2",x"87",x"f7"),
  1088 => (x"78",x"c0",x"48",x"e8"),
  1089 => (x"e0",x"c0",x"49",x"c1"),
  1090 => (x"fb",x"26",x"87",x"ff"),
  1091 => (x"6f",x"4c",x"87",x"dd"),
  1092 => (x"6e",x"69",x"64",x"61"),
  1093 => (x"2e",x"2e",x"2e",x"67"),
  1094 => (x"5b",x"5e",x"0e",x"00"),
  1095 => (x"4b",x"71",x"0e",x"5c"),
  1096 => (x"c0",x"f4",x"c2",x"4a"),
  1097 => (x"49",x"72",x"82",x"bf"),
  1098 => (x"70",x"87",x"c8",x"fb"),
  1099 => (x"c4",x"02",x"9c",x"4c"),
  1100 => (x"dd",x"e5",x"49",x"87"),
  1101 => (x"c0",x"f4",x"c2",x"87"),
  1102 => (x"c1",x"78",x"c0",x"48"),
  1103 => (x"c8",x"e0",x"c0",x"49"),
  1104 => (x"87",x"e9",x"fa",x"87"),
  1105 => (x"5c",x"5b",x"5e",x"0e"),
  1106 => (x"86",x"f4",x"0e",x"5d"),
  1107 => (x"4d",x"f6",x"e6",x"c2"),
  1108 => (x"a6",x"c4",x"4c",x"c0"),
  1109 => (x"c2",x"78",x"c0",x"48"),
  1110 => (x"49",x"bf",x"c0",x"f4"),
  1111 => (x"c1",x"06",x"a9",x"c0"),
  1112 => (x"e6",x"c2",x"87",x"c1"),
  1113 => (x"02",x"98",x"48",x"f6"),
  1114 => (x"c0",x"87",x"f8",x"c0"),
  1115 => (x"c8",x"1e",x"d5",x"f7"),
  1116 => (x"87",x"c7",x"02",x"66"),
  1117 => (x"c0",x"48",x"a6",x"c4"),
  1118 => (x"c4",x"87",x"c5",x"78"),
  1119 => (x"78",x"c1",x"48",x"a6"),
  1120 => (x"e5",x"49",x"66",x"c4"),
  1121 => (x"86",x"c4",x"87",x"c4"),
  1122 => (x"84",x"c1",x"4d",x"70"),
  1123 => (x"c1",x"48",x"66",x"c4"),
  1124 => (x"58",x"a6",x"c8",x"80"),
  1125 => (x"bf",x"c0",x"f4",x"c2"),
  1126 => (x"c6",x"03",x"ac",x"49"),
  1127 => (x"05",x"9d",x"75",x"87"),
  1128 => (x"c0",x"87",x"c8",x"ff"),
  1129 => (x"02",x"9d",x"75",x"4c"),
  1130 => (x"c0",x"87",x"e0",x"c3"),
  1131 => (x"c8",x"1e",x"d5",x"f7"),
  1132 => (x"87",x"c7",x"02",x"66"),
  1133 => (x"c0",x"48",x"a6",x"cc"),
  1134 => (x"cc",x"87",x"c5",x"78"),
  1135 => (x"78",x"c1",x"48",x"a6"),
  1136 => (x"e4",x"49",x"66",x"cc"),
  1137 => (x"86",x"c4",x"87",x"c4"),
  1138 => (x"98",x"48",x"7e",x"70"),
  1139 => (x"87",x"e8",x"c2",x"02"),
  1140 => (x"97",x"81",x"cb",x"49"),
  1141 => (x"99",x"d0",x"49",x"69"),
  1142 => (x"87",x"d6",x"c1",x"02"),
  1143 => (x"4a",x"d9",x"c4",x"c1"),
  1144 => (x"91",x"cb",x"49",x"74"),
  1145 => (x"81",x"ef",x"e9",x"c1"),
  1146 => (x"81",x"c8",x"79",x"72"),
  1147 => (x"74",x"51",x"ff",x"c3"),
  1148 => (x"c2",x"91",x"de",x"49"),
  1149 => (x"71",x"4d",x"d4",x"f4"),
  1150 => (x"97",x"c1",x"c2",x"85"),
  1151 => (x"49",x"a5",x"c1",x"7d"),
  1152 => (x"c2",x"51",x"e0",x"c0"),
  1153 => (x"bf",x"97",x"c6",x"ef"),
  1154 => (x"c1",x"87",x"d2",x"02"),
  1155 => (x"4b",x"a5",x"c2",x"84"),
  1156 => (x"4a",x"c6",x"ef",x"c2"),
  1157 => (x"fa",x"fe",x"49",x"db"),
  1158 => (x"db",x"c1",x"87",x"cd"),
  1159 => (x"49",x"a5",x"cd",x"87"),
  1160 => (x"84",x"c1",x"51",x"c0"),
  1161 => (x"6e",x"4b",x"a5",x"c2"),
  1162 => (x"fe",x"49",x"cb",x"4a"),
  1163 => (x"c1",x"87",x"f8",x"f9"),
  1164 => (x"c2",x"c1",x"87",x"c6"),
  1165 => (x"49",x"74",x"4a",x"d4"),
  1166 => (x"e9",x"c1",x"91",x"cb"),
  1167 => (x"79",x"72",x"81",x"ef"),
  1168 => (x"97",x"c6",x"ef",x"c2"),
  1169 => (x"87",x"d8",x"02",x"bf"),
  1170 => (x"91",x"de",x"49",x"74"),
  1171 => (x"f4",x"c2",x"84",x"c1"),
  1172 => (x"83",x"71",x"4b",x"d4"),
  1173 => (x"4a",x"c6",x"ef",x"c2"),
  1174 => (x"f9",x"fe",x"49",x"dd"),
  1175 => (x"87",x"d8",x"87",x"c9"),
  1176 => (x"93",x"de",x"4b",x"74"),
  1177 => (x"83",x"d4",x"f4",x"c2"),
  1178 => (x"c0",x"49",x"a3",x"cb"),
  1179 => (x"73",x"84",x"c1",x"51"),
  1180 => (x"49",x"cb",x"4a",x"6e"),
  1181 => (x"87",x"ef",x"f8",x"fe"),
  1182 => (x"c1",x"48",x"66",x"c4"),
  1183 => (x"58",x"a6",x"c8",x"80"),
  1184 => (x"c0",x"03",x"ac",x"c7"),
  1185 => (x"05",x"6e",x"87",x"c5"),
  1186 => (x"74",x"87",x"e0",x"fc"),
  1187 => (x"f5",x"8e",x"f4",x"48"),
  1188 => (x"73",x"1e",x"87",x"d9"),
  1189 => (x"49",x"4b",x"71",x"1e"),
  1190 => (x"e9",x"c1",x"91",x"cb"),
  1191 => (x"a1",x"c8",x"81",x"ef"),
  1192 => (x"f8",x"e8",x"c1",x"4a"),
  1193 => (x"c9",x"50",x"12",x"48"),
  1194 => (x"fa",x"c0",x"4a",x"a1"),
  1195 => (x"50",x"12",x"48",x"fc"),
  1196 => (x"e8",x"c1",x"81",x"ca"),
  1197 => (x"50",x"11",x"48",x"f9"),
  1198 => (x"97",x"f9",x"e8",x"c1"),
  1199 => (x"c0",x"1e",x"49",x"bf"),
  1200 => (x"87",x"ee",x"f5",x"49"),
  1201 => (x"48",x"e8",x"f3",x"c2"),
  1202 => (x"49",x"c1",x"78",x"de"),
  1203 => (x"26",x"87",x"fa",x"d9"),
  1204 => (x"1e",x"87",x"dc",x"f4"),
  1205 => (x"cb",x"49",x"4a",x"71"),
  1206 => (x"ef",x"e9",x"c1",x"91"),
  1207 => (x"11",x"81",x"c8",x"81"),
  1208 => (x"ec",x"f3",x"c2",x"48"),
  1209 => (x"c0",x"f4",x"c2",x"58"),
  1210 => (x"c1",x"78",x"c0",x"48"),
  1211 => (x"87",x"d9",x"d9",x"49"),
  1212 => (x"c0",x"1e",x"4f",x"26"),
  1213 => (x"fc",x"fe",x"c0",x"49"),
  1214 => (x"1e",x"4f",x"26",x"87"),
  1215 => (x"d2",x"02",x"99",x"71"),
  1216 => (x"c4",x"eb",x"c1",x"87"),
  1217 => (x"f7",x"50",x"c0",x"48"),
  1218 => (x"d3",x"cb",x"c1",x"80"),
  1219 => (x"dd",x"e9",x"c1",x"40"),
  1220 => (x"c1",x"87",x"ce",x"78"),
  1221 => (x"c1",x"48",x"c0",x"eb"),
  1222 => (x"fc",x"78",x"fe",x"e8"),
  1223 => (x"f2",x"cb",x"c1",x"80"),
  1224 => (x"0e",x"4f",x"26",x"78"),
  1225 => (x"5d",x"5c",x"5b",x"5e"),
  1226 => (x"71",x"86",x"f4",x"0e"),
  1227 => (x"91",x"cb",x"49",x"4d"),
  1228 => (x"81",x"ef",x"e9",x"c1"),
  1229 => (x"ca",x"4a",x"a1",x"c8"),
  1230 => (x"a6",x"c4",x"7e",x"a1"),
  1231 => (x"f0",x"f7",x"c2",x"48"),
  1232 => (x"97",x"6e",x"78",x"bf"),
  1233 => (x"66",x"c4",x"4b",x"bf"),
  1234 => (x"70",x"28",x"73",x"48"),
  1235 => (x"48",x"12",x"4c",x"4b"),
  1236 => (x"70",x"58",x"a6",x"cc"),
  1237 => (x"c9",x"84",x"c1",x"9c"),
  1238 => (x"49",x"69",x"97",x"81"),
  1239 => (x"c2",x"04",x"ac",x"b7"),
  1240 => (x"6e",x"4c",x"c0",x"87"),
  1241 => (x"c8",x"4a",x"bf",x"97"),
  1242 => (x"31",x"72",x"49",x"66"),
  1243 => (x"66",x"c4",x"b9",x"ff"),
  1244 => (x"72",x"48",x"74",x"99"),
  1245 => (x"48",x"4a",x"70",x"30"),
  1246 => (x"f7",x"c2",x"b0",x"71"),
  1247 => (x"e9",x"c0",x"58",x"f4"),
  1248 => (x"49",x"c0",x"87",x"ce"),
  1249 => (x"75",x"87",x"c2",x"d7"),
  1250 => (x"c3",x"fb",x"c0",x"49"),
  1251 => (x"f1",x"8e",x"f4",x"87"),
  1252 => (x"73",x"1e",x"87",x"d9"),
  1253 => (x"49",x"4b",x"71",x"1e"),
  1254 => (x"73",x"87",x"c8",x"fe"),
  1255 => (x"87",x"c3",x"fe",x"49"),
  1256 => (x"1e",x"87",x"cc",x"f1"),
  1257 => (x"4b",x"71",x"1e",x"73"),
  1258 => (x"02",x"4a",x"a3",x"c6"),
  1259 => (x"8a",x"c1",x"87",x"dc"),
  1260 => (x"87",x"e4",x"c0",x"02"),
  1261 => (x"e8",x"c1",x"02",x"8a"),
  1262 => (x"c1",x"02",x"8a",x"87"),
  1263 => (x"02",x"8a",x"87",x"ca"),
  1264 => (x"8a",x"87",x"ef",x"c0"),
  1265 => (x"c1",x"87",x"d9",x"02"),
  1266 => (x"f3",x"c2",x"87",x"e9"),
  1267 => (x"78",x"df",x"48",x"e8"),
  1268 => (x"f4",x"d5",x"49",x"c1"),
  1269 => (x"87",x"e6",x"c1",x"87"),
  1270 => (x"f6",x"fb",x"49",x"c7"),
  1271 => (x"87",x"de",x"c1",x"87"),
  1272 => (x"bf",x"c0",x"f4",x"c2"),
  1273 => (x"87",x"cb",x"c1",x"02"),
  1274 => (x"c2",x"88",x"c1",x"48"),
  1275 => (x"c1",x"58",x"c4",x"f4"),
  1276 => (x"f4",x"c2",x"87",x"c1"),
  1277 => (x"c0",x"02",x"bf",x"c4"),
  1278 => (x"f4",x"c2",x"87",x"f9"),
  1279 => (x"c1",x"48",x"bf",x"c0"),
  1280 => (x"c4",x"f4",x"c2",x"80"),
  1281 => (x"87",x"eb",x"c0",x"58"),
  1282 => (x"bf",x"c0",x"f4",x"c2"),
  1283 => (x"c2",x"89",x"c6",x"49"),
  1284 => (x"c0",x"59",x"c4",x"f4"),
  1285 => (x"da",x"03",x"a9",x"b7"),
  1286 => (x"c0",x"f4",x"c2",x"87"),
  1287 => (x"d2",x"78",x"c0",x"48"),
  1288 => (x"c4",x"f4",x"c2",x"87"),
  1289 => (x"87",x"cb",x"02",x"bf"),
  1290 => (x"bf",x"c0",x"f4",x"c2"),
  1291 => (x"c2",x"80",x"c6",x"48"),
  1292 => (x"c0",x"58",x"c4",x"f4"),
  1293 => (x"87",x"d1",x"d4",x"49"),
  1294 => (x"f8",x"c0",x"49",x"73"),
  1295 => (x"ee",x"ee",x"87",x"d2"),
  1296 => (x"5b",x"5e",x"0e",x"87"),
  1297 => (x"ff",x"0e",x"5d",x"5c"),
  1298 => (x"a6",x"dc",x"86",x"d0"),
  1299 => (x"cc",x"4d",x"c0",x"59"),
  1300 => (x"c4",x"c1",x"48",x"a6"),
  1301 => (x"80",x"c4",x"78",x"66"),
  1302 => (x"80",x"c4",x"78",x"c1"),
  1303 => (x"f4",x"c2",x"78",x"c1"),
  1304 => (x"78",x"c1",x"48",x"c4"),
  1305 => (x"bf",x"e8",x"f3",x"c2"),
  1306 => (x"de",x"48",x"6e",x"7e"),
  1307 => (x"87",x"c9",x"05",x"a8"),
  1308 => (x"70",x"87",x"d1",x"f3"),
  1309 => (x"f9",x"d1",x"4d",x"49"),
  1310 => (x"df",x"48",x"6e",x"87"),
  1311 => (x"eb",x"c1",x"05",x"a8"),
  1312 => (x"66",x"c0",x"c1",x"87"),
  1313 => (x"69",x"81",x"c4",x"49"),
  1314 => (x"dd",x"e4",x"c1",x"7e"),
  1315 => (x"d0",x"49",x"6e",x"48"),
  1316 => (x"41",x"20",x"4a",x"a1"),
  1317 => (x"f9",x"05",x"aa",x"71"),
  1318 => (x"d2",x"ca",x"c1",x"87"),
  1319 => (x"66",x"c0",x"c1",x"4a"),
  1320 => (x"c1",x"0a",x"7a",x"0a"),
  1321 => (x"c9",x"49",x"66",x"c0"),
  1322 => (x"c1",x"51",x"df",x"81"),
  1323 => (x"ca",x"49",x"66",x"c0"),
  1324 => (x"51",x"d3",x"c1",x"81"),
  1325 => (x"49",x"66",x"c0",x"c1"),
  1326 => (x"a1",x"c4",x"81",x"cb"),
  1327 => (x"48",x"a6",x"c4",x"4b"),
  1328 => (x"1e",x"71",x"78",x"6b"),
  1329 => (x"e4",x"c1",x"1e",x"72"),
  1330 => (x"66",x"cc",x"48",x"ed"),
  1331 => (x"4a",x"a1",x"d0",x"49"),
  1332 => (x"aa",x"71",x"41",x"20"),
  1333 => (x"26",x"87",x"f9",x"05"),
  1334 => (x"72",x"49",x"26",x"4a"),
  1335 => (x"4a",x"a1",x"c9",x"79"),
  1336 => (x"81",x"ca",x"52",x"df"),
  1337 => (x"c2",x"51",x"d4",x"c1"),
  1338 => (x"87",x"c6",x"d0",x"4d"),
  1339 => (x"87",x"de",x"df",x"ff"),
  1340 => (x"ff",x"87",x"c0",x"e0"),
  1341 => (x"70",x"87",x"cc",x"df"),
  1342 => (x"ac",x"fb",x"c0",x"4c"),
  1343 => (x"87",x"fa",x"c1",x"02"),
  1344 => (x"c1",x"05",x"66",x"d8"),
  1345 => (x"c0",x"c1",x"87",x"eb"),
  1346 => (x"82",x"c4",x"4a",x"66"),
  1347 => (x"1e",x"72",x"7e",x"6a"),
  1348 => (x"48",x"fd",x"e4",x"c1"),
  1349 => (x"c8",x"49",x"66",x"c4"),
  1350 => (x"41",x"20",x"4a",x"a1"),
  1351 => (x"f9",x"05",x"aa",x"71"),
  1352 => (x"26",x"51",x"10",x"87"),
  1353 => (x"66",x"c0",x"c1",x"4a"),
  1354 => (x"d2",x"ca",x"c1",x"48"),
  1355 => (x"c7",x"49",x"6a",x"78"),
  1356 => (x"c1",x"51",x"74",x"81"),
  1357 => (x"c8",x"49",x"66",x"c0"),
  1358 => (x"c1",x"51",x"c1",x"81"),
  1359 => (x"c9",x"49",x"66",x"c0"),
  1360 => (x"c1",x"51",x"c0",x"81"),
  1361 => (x"ca",x"49",x"66",x"c0"),
  1362 => (x"c1",x"51",x"c0",x"81"),
  1363 => (x"6a",x"1e",x"d8",x"1e"),
  1364 => (x"ff",x"81",x"c8",x"49"),
  1365 => (x"c8",x"87",x"f0",x"de"),
  1366 => (x"66",x"c4",x"c1",x"86"),
  1367 => (x"01",x"a8",x"c0",x"48"),
  1368 => (x"4d",x"c1",x"87",x"c4"),
  1369 => (x"c4",x"c1",x"87",x"cf"),
  1370 => (x"88",x"c1",x"48",x"66"),
  1371 => (x"c4",x"58",x"a6",x"d0"),
  1372 => (x"fe",x"dd",x"ff",x"87"),
  1373 => (x"48",x"a6",x"d0",x"87"),
  1374 => (x"a6",x"cc",x"78",x"c2"),
  1375 => (x"02",x"9c",x"74",x"5d"),
  1376 => (x"cc",x"87",x"e8",x"cd"),
  1377 => (x"c8",x"c1",x"5d",x"a6"),
  1378 => (x"cd",x"03",x"ad",x"66"),
  1379 => (x"a6",x"dc",x"87",x"dd"),
  1380 => (x"e8",x"78",x"c0",x"48"),
  1381 => (x"ff",x"78",x"c0",x"80"),
  1382 => (x"70",x"87",x"e8",x"dc"),
  1383 => (x"ac",x"d0",x"c1",x"4c"),
  1384 => (x"87",x"db",x"c2",x"05"),
  1385 => (x"ff",x"7e",x"66",x"c4"),
  1386 => (x"70",x"87",x"cb",x"df"),
  1387 => (x"59",x"a6",x"c8",x"49"),
  1388 => (x"87",x"cf",x"dc",x"ff"),
  1389 => (x"ec",x"c0",x"4c",x"70"),
  1390 => (x"ed",x"c1",x"05",x"ac"),
  1391 => (x"49",x"66",x"c8",x"87"),
  1392 => (x"c0",x"c1",x"91",x"cb"),
  1393 => (x"a1",x"c4",x"81",x"66"),
  1394 => (x"c8",x"4d",x"6a",x"4a"),
  1395 => (x"66",x"c4",x"4a",x"a1"),
  1396 => (x"d3",x"cb",x"c1",x"52"),
  1397 => (x"ea",x"db",x"ff",x"79"),
  1398 => (x"9c",x"4c",x"70",x"87"),
  1399 => (x"c0",x"87",x"d9",x"02"),
  1400 => (x"d3",x"02",x"ac",x"fb"),
  1401 => (x"ff",x"55",x"74",x"87"),
  1402 => (x"70",x"87",x"d8",x"db"),
  1403 => (x"c7",x"02",x"9c",x"4c"),
  1404 => (x"ac",x"fb",x"c0",x"87"),
  1405 => (x"87",x"ed",x"ff",x"05"),
  1406 => (x"c2",x"55",x"e0",x"c0"),
  1407 => (x"97",x"c0",x"55",x"c1"),
  1408 => (x"49",x"66",x"d8",x"7d"),
  1409 => (x"db",x"05",x"a9",x"6e"),
  1410 => (x"48",x"66",x"c8",x"87"),
  1411 => (x"04",x"a8",x"66",x"cc"),
  1412 => (x"66",x"c8",x"87",x"ca"),
  1413 => (x"cc",x"80",x"c1",x"48"),
  1414 => (x"87",x"c8",x"58",x"a6"),
  1415 => (x"c1",x"48",x"66",x"cc"),
  1416 => (x"58",x"a6",x"d0",x"88"),
  1417 => (x"87",x"db",x"da",x"ff"),
  1418 => (x"d0",x"c1",x"4c",x"70"),
  1419 => (x"87",x"c8",x"05",x"ac"),
  1420 => (x"c1",x"48",x"66",x"d4"),
  1421 => (x"58",x"a6",x"d8",x"80"),
  1422 => (x"02",x"ac",x"d0",x"c1"),
  1423 => (x"c0",x"87",x"e5",x"fd"),
  1424 => (x"d8",x"48",x"a6",x"e0"),
  1425 => (x"66",x"c4",x"78",x"66"),
  1426 => (x"66",x"e0",x"c0",x"48"),
  1427 => (x"ec",x"c9",x"05",x"a8"),
  1428 => (x"a6",x"e4",x"c0",x"87"),
  1429 => (x"74",x"78",x"c0",x"48"),
  1430 => (x"88",x"fb",x"c0",x"48"),
  1431 => (x"98",x"48",x"7e",x"70"),
  1432 => (x"87",x"ee",x"c9",x"02"),
  1433 => (x"70",x"88",x"cb",x"48"),
  1434 => (x"02",x"98",x"48",x"7e"),
  1435 => (x"48",x"87",x"ce",x"c1"),
  1436 => (x"7e",x"70",x"88",x"c9"),
  1437 => (x"c4",x"02",x"98",x"48"),
  1438 => (x"c4",x"48",x"87",x"c2"),
  1439 => (x"48",x"7e",x"70",x"88"),
  1440 => (x"87",x"ce",x"02",x"98"),
  1441 => (x"70",x"88",x"c1",x"48"),
  1442 => (x"02",x"98",x"48",x"7e"),
  1443 => (x"c8",x"87",x"ed",x"c3"),
  1444 => (x"a6",x"dc",x"87",x"e2"),
  1445 => (x"78",x"f0",x"c0",x"48"),
  1446 => (x"87",x"e7",x"d8",x"ff"),
  1447 => (x"ec",x"c0",x"4c",x"70"),
  1448 => (x"c4",x"c0",x"02",x"ac"),
  1449 => (x"a6",x"e0",x"c0",x"87"),
  1450 => (x"ac",x"ec",x"c0",x"5c"),
  1451 => (x"87",x"cd",x"c0",x"02"),
  1452 => (x"87",x"cf",x"d8",x"ff"),
  1453 => (x"ec",x"c0",x"4c",x"70"),
  1454 => (x"f3",x"ff",x"05",x"ac"),
  1455 => (x"ac",x"ec",x"c0",x"87"),
  1456 => (x"87",x"c4",x"c0",x"02"),
  1457 => (x"87",x"fb",x"d7",x"ff"),
  1458 => (x"1e",x"ca",x"1e",x"c0"),
  1459 => (x"cb",x"49",x"66",x"d0"),
  1460 => (x"66",x"c8",x"c1",x"91"),
  1461 => (x"cc",x"80",x"71",x"48"),
  1462 => (x"66",x"c8",x"58",x"a6"),
  1463 => (x"d0",x"80",x"c4",x"48"),
  1464 => (x"66",x"cc",x"58",x"a6"),
  1465 => (x"d8",x"ff",x"49",x"bf"),
  1466 => (x"1e",x"c1",x"87",x"dd"),
  1467 => (x"66",x"d4",x"1e",x"de"),
  1468 => (x"d8",x"ff",x"49",x"bf"),
  1469 => (x"86",x"d0",x"87",x"d1"),
  1470 => (x"09",x"c0",x"49",x"70"),
  1471 => (x"a6",x"ec",x"c0",x"89"),
  1472 => (x"66",x"e8",x"c0",x"59"),
  1473 => (x"06",x"a8",x"c0",x"48"),
  1474 => (x"c0",x"87",x"ee",x"c0"),
  1475 => (x"dd",x"48",x"66",x"e8"),
  1476 => (x"e4",x"c0",x"03",x"a8"),
  1477 => (x"bf",x"66",x"c4",x"87"),
  1478 => (x"66",x"e8",x"c0",x"49"),
  1479 => (x"51",x"e0",x"c0",x"81"),
  1480 => (x"49",x"66",x"e8",x"c0"),
  1481 => (x"66",x"c4",x"81",x"c1"),
  1482 => (x"c1",x"c2",x"81",x"bf"),
  1483 => (x"66",x"e8",x"c0",x"51"),
  1484 => (x"c4",x"81",x"c2",x"49"),
  1485 => (x"c0",x"81",x"bf",x"66"),
  1486 => (x"c1",x"48",x"6e",x"51"),
  1487 => (x"6e",x"78",x"d2",x"ca"),
  1488 => (x"d0",x"81",x"c8",x"49"),
  1489 => (x"49",x"6e",x"51",x"66"),
  1490 => (x"66",x"d4",x"81",x"c9"),
  1491 => (x"ca",x"49",x"6e",x"51"),
  1492 => (x"51",x"66",x"dc",x"81"),
  1493 => (x"c1",x"48",x"66",x"d0"),
  1494 => (x"58",x"a6",x"d4",x"80"),
  1495 => (x"cc",x"48",x"66",x"c8"),
  1496 => (x"c0",x"04",x"a8",x"66"),
  1497 => (x"66",x"c8",x"87",x"cb"),
  1498 => (x"cc",x"80",x"c1",x"48"),
  1499 => (x"e1",x"c5",x"58",x"a6"),
  1500 => (x"48",x"66",x"cc",x"87"),
  1501 => (x"a6",x"d0",x"88",x"c1"),
  1502 => (x"87",x"d6",x"c5",x"58"),
  1503 => (x"87",x"f6",x"d7",x"ff"),
  1504 => (x"ec",x"c0",x"49",x"70"),
  1505 => (x"d7",x"ff",x"59",x"a6"),
  1506 => (x"49",x"70",x"87",x"ec"),
  1507 => (x"59",x"a6",x"e0",x"c0"),
  1508 => (x"c0",x"48",x"66",x"dc"),
  1509 => (x"c0",x"05",x"a8",x"ec"),
  1510 => (x"a6",x"dc",x"87",x"ca"),
  1511 => (x"66",x"e8",x"c0",x"48"),
  1512 => (x"87",x"c4",x"c0",x"78"),
  1513 => (x"87",x"db",x"d4",x"ff"),
  1514 => (x"cb",x"49",x"66",x"c8"),
  1515 => (x"66",x"c0",x"c1",x"91"),
  1516 => (x"70",x"80",x"71",x"48"),
  1517 => (x"82",x"c8",x"4a",x"7e"),
  1518 => (x"81",x"ca",x"49",x"6e"),
  1519 => (x"51",x"66",x"e8",x"c0"),
  1520 => (x"c1",x"49",x"66",x"dc"),
  1521 => (x"66",x"e8",x"c0",x"81"),
  1522 => (x"71",x"48",x"c1",x"89"),
  1523 => (x"c1",x"49",x"70",x"30"),
  1524 => (x"7a",x"97",x"71",x"89"),
  1525 => (x"bf",x"f0",x"f7",x"c2"),
  1526 => (x"66",x"e8",x"c0",x"49"),
  1527 => (x"4a",x"6a",x"97",x"29"),
  1528 => (x"c0",x"98",x"71",x"48"),
  1529 => (x"6e",x"58",x"a6",x"f0"),
  1530 => (x"69",x"81",x"c4",x"49"),
  1531 => (x"66",x"e0",x"c0",x"4d"),
  1532 => (x"a8",x"66",x"c4",x"48"),
  1533 => (x"87",x"c8",x"c0",x"02"),
  1534 => (x"c0",x"48",x"a6",x"c4"),
  1535 => (x"87",x"c5",x"c0",x"78"),
  1536 => (x"c1",x"48",x"a6",x"c4"),
  1537 => (x"1e",x"66",x"c4",x"78"),
  1538 => (x"75",x"1e",x"e0",x"c0"),
  1539 => (x"f6",x"d3",x"ff",x"49"),
  1540 => (x"70",x"86",x"c8",x"87"),
  1541 => (x"ac",x"b7",x"c0",x"4c"),
  1542 => (x"87",x"d4",x"c1",x"06"),
  1543 => (x"e0",x"c0",x"85",x"74"),
  1544 => (x"75",x"89",x"74",x"49"),
  1545 => (x"c6",x"e5",x"c1",x"4b"),
  1546 => (x"e1",x"fe",x"71",x"4a"),
  1547 => (x"85",x"c2",x"87",x"f9"),
  1548 => (x"48",x"66",x"e4",x"c0"),
  1549 => (x"e8",x"c0",x"80",x"c1"),
  1550 => (x"ec",x"c0",x"58",x"a6"),
  1551 => (x"81",x"c1",x"49",x"66"),
  1552 => (x"c0",x"02",x"a9",x"70"),
  1553 => (x"a6",x"c4",x"87",x"c8"),
  1554 => (x"c0",x"78",x"c0",x"48"),
  1555 => (x"a6",x"c4",x"87",x"c5"),
  1556 => (x"c4",x"78",x"c1",x"48"),
  1557 => (x"a4",x"c2",x"1e",x"66"),
  1558 => (x"48",x"e0",x"c0",x"49"),
  1559 => (x"49",x"70",x"88",x"71"),
  1560 => (x"ff",x"49",x"75",x"1e"),
  1561 => (x"c8",x"87",x"e0",x"d2"),
  1562 => (x"a8",x"b7",x"c0",x"86"),
  1563 => (x"87",x"c0",x"ff",x"01"),
  1564 => (x"02",x"66",x"e4",x"c0"),
  1565 => (x"6e",x"87",x"d1",x"c0"),
  1566 => (x"c0",x"81",x"c9",x"49"),
  1567 => (x"6e",x"51",x"66",x"e4"),
  1568 => (x"e3",x"cc",x"c1",x"48"),
  1569 => (x"87",x"cc",x"c0",x"78"),
  1570 => (x"81",x"c9",x"49",x"6e"),
  1571 => (x"48",x"6e",x"51",x"c2"),
  1572 => (x"78",x"d2",x"ce",x"c1"),
  1573 => (x"cc",x"48",x"66",x"c8"),
  1574 => (x"c0",x"04",x"a8",x"66"),
  1575 => (x"66",x"c8",x"87",x"cb"),
  1576 => (x"cc",x"80",x"c1",x"48"),
  1577 => (x"e9",x"c0",x"58",x"a6"),
  1578 => (x"48",x"66",x"cc",x"87"),
  1579 => (x"a6",x"d0",x"88",x"c1"),
  1580 => (x"87",x"de",x"c0",x"58"),
  1581 => (x"87",x"fb",x"d0",x"ff"),
  1582 => (x"d5",x"c0",x"4c",x"70"),
  1583 => (x"ac",x"c6",x"c1",x"87"),
  1584 => (x"87",x"c8",x"c0",x"05"),
  1585 => (x"c1",x"48",x"66",x"d0"),
  1586 => (x"58",x"a6",x"d4",x"80"),
  1587 => (x"87",x"e3",x"d0",x"ff"),
  1588 => (x"66",x"d4",x"4c",x"70"),
  1589 => (x"d8",x"80",x"c1",x"48"),
  1590 => (x"9c",x"74",x"58",x"a6"),
  1591 => (x"87",x"cb",x"c0",x"02"),
  1592 => (x"c1",x"48",x"66",x"c8"),
  1593 => (x"04",x"a8",x"66",x"c8"),
  1594 => (x"c8",x"87",x"e3",x"f2"),
  1595 => (x"cf",x"ff",x"4d",x"66"),
  1596 => (x"ad",x"c7",x"87",x"f8"),
  1597 => (x"87",x"de",x"c0",x"03"),
  1598 => (x"48",x"c4",x"f4",x"c2"),
  1599 => (x"49",x"75",x"78",x"c0"),
  1600 => (x"c0",x"c1",x"91",x"cb"),
  1601 => (x"a1",x"c4",x"81",x"66"),
  1602 => (x"c0",x"4a",x"6a",x"4a"),
  1603 => (x"85",x"c1",x"79",x"52"),
  1604 => (x"ff",x"04",x"ad",x"c7"),
  1605 => (x"d0",x"ff",x"87",x"e2"),
  1606 => (x"ce",x"db",x"ff",x"8e"),
  1607 => (x"61",x"6f",x"4c",x"87"),
  1608 => (x"65",x"53",x"20",x"64"),
  1609 => (x"6e",x"69",x"74",x"74"),
  1610 => (x"81",x"20",x"73",x"67"),
  1611 => (x"76",x"61",x"53",x"00"),
  1612 => (x"65",x"53",x"20",x"65"),
  1613 => (x"6e",x"69",x"74",x"74"),
  1614 => (x"81",x"20",x"73",x"67"),
  1615 => (x"61",x"6f",x"4c",x"00"),
  1616 => (x"2e",x"2a",x"20",x"64"),
  1617 => (x"20",x"3a",x"00",x"20"),
  1618 => (x"1e",x"73",x"1e",x"00"),
  1619 => (x"02",x"9b",x"4b",x"71"),
  1620 => (x"f4",x"c2",x"87",x"c6"),
  1621 => (x"78",x"c0",x"48",x"c0"),
  1622 => (x"f4",x"c2",x"1e",x"c7"),
  1623 => (x"1e",x"49",x"bf",x"c0"),
  1624 => (x"1e",x"ef",x"e9",x"c1"),
  1625 => (x"bf",x"e8",x"f3",x"c2"),
  1626 => (x"87",x"d5",x"eb",x"49"),
  1627 => (x"f3",x"c2",x"86",x"cc"),
  1628 => (x"e6",x"49",x"bf",x"e8"),
  1629 => (x"9b",x"73",x"87",x"c5"),
  1630 => (x"c1",x"87",x"c8",x"02"),
  1631 => (x"c0",x"49",x"ef",x"e9"),
  1632 => (x"ff",x"87",x"df",x"e4"),
  1633 => (x"1e",x"87",x"e8",x"d9"),
  1634 => (x"49",x"e3",x"e6",x"c1"),
  1635 => (x"87",x"cc",x"fe",x"c0"),
  1636 => (x"48",x"f8",x"e8",x"c1"),
  1637 => (x"eb",x"c1",x"50",x"c0"),
  1638 => (x"ff",x"49",x"bf",x"d2"),
  1639 => (x"c0",x"87",x"de",x"d4"),
  1640 => (x"4f",x"4f",x"26",x"48"),
  1641 => (x"20",x"43",x"49",x"52"),
  1642 => (x"43",x"20",x"20",x"20"),
  1643 => (x"1e",x"00",x"47",x"46"),
  1644 => (x"c1",x"87",x"c6",x"c8"),
  1645 => (x"87",x"d1",x"fe",x"49"),
  1646 => (x"87",x"d3",x"e4",x"fe"),
  1647 => (x"cd",x"02",x"98",x"70"),
  1648 => (x"ce",x"ed",x"fe",x"87"),
  1649 => (x"02",x"98",x"70",x"87"),
  1650 => (x"4a",x"c1",x"87",x"c4"),
  1651 => (x"4a",x"c0",x"87",x"c2"),
  1652 => (x"ce",x"05",x"9a",x"72"),
  1653 => (x"c1",x"1e",x"c0",x"87"),
  1654 => (x"c0",x"49",x"ff",x"e7"),
  1655 => (x"c4",x"87",x"e9",x"f2"),
  1656 => (x"c0",x"87",x"fe",x"86"),
  1657 => (x"ca",x"e8",x"c1",x"1e"),
  1658 => (x"db",x"f2",x"c0",x"49"),
  1659 => (x"fe",x"1e",x"c0",x"87"),
  1660 => (x"49",x"70",x"87",x"d5"),
  1661 => (x"87",x"d0",x"f2",x"c0"),
  1662 => (x"f8",x"87",x"fd",x"c3"),
  1663 => (x"53",x"4f",x"26",x"8e"),
  1664 => (x"61",x"66",x"20",x"44"),
  1665 => (x"64",x"65",x"6c",x"69"),
  1666 => (x"6f",x"42",x"00",x"2e"),
  1667 => (x"6e",x"69",x"74",x"6f"),
  1668 => (x"2e",x"2e",x"2e",x"67"),
  1669 => (x"e7",x"c0",x"1e",x"00"),
  1670 => (x"f5",x"c0",x"87",x"cd"),
  1671 => (x"87",x"f6",x"87",x"f9"),
  1672 => (x"c2",x"1e",x"4f",x"26"),
  1673 => (x"c0",x"48",x"c0",x"f4"),
  1674 => (x"e8",x"f3",x"c2",x"78"),
  1675 => (x"fd",x"78",x"c0",x"48"),
  1676 => (x"87",x"e1",x"87",x"fd"),
  1677 => (x"4f",x"26",x"48",x"c0"),
  1678 => (x"00",x"01",x"00",x"00"),
  1679 => (x"20",x"20",x"00",x"00"),
  1680 => (x"20",x"20",x"20",x"20"),
  1681 => (x"20",x"20",x"20",x"20"),
  1682 => (x"45",x"20",x"20",x"20"),
  1683 => (x"20",x"74",x"69",x"78"),
  1684 => (x"20",x"20",x"20",x"20"),
  1685 => (x"20",x"20",x"20",x"20"),
  1686 => (x"81",x"20",x"20",x"20"),
  1687 => (x"20",x"20",x"80",x"00"),
  1688 => (x"20",x"20",x"20",x"20"),
  1689 => (x"20",x"20",x"20",x"20"),
  1690 => (x"61",x"42",x"20",x"20"),
  1691 => (x"94",x"00",x"6b",x"63"),
  1692 => (x"14",x"00",x"00",x"10"),
  1693 => (x"00",x"00",x"00",x"2d"),
  1694 => (x"10",x"94",x"00",x"00"),
  1695 => (x"2d",x"32",x"00",x"00"),
  1696 => (x"00",x"00",x"00",x"00"),
  1697 => (x"00",x"10",x"94",x"00"),
  1698 => (x"00",x"2d",x"50",x"00"),
  1699 => (x"00",x"00",x"00",x"00"),
  1700 => (x"00",x"00",x"10",x"94"),
  1701 => (x"00",x"00",x"2d",x"6e"),
  1702 => (x"94",x"00",x"00",x"00"),
  1703 => (x"8c",x"00",x"00",x"10"),
  1704 => (x"00",x"00",x"00",x"2d"),
  1705 => (x"10",x"94",x"00",x"00"),
  1706 => (x"2d",x"aa",x"00",x"00"),
  1707 => (x"00",x"00",x"00",x"00"),
  1708 => (x"00",x"10",x"94",x"00"),
  1709 => (x"00",x"2d",x"c8",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"12",x"d3"),
  1712 => (x"00",x"00",x"00",x"00"),
  1713 => (x"a3",x"00",x"00",x"00"),
  1714 => (x"00",x"00",x"00",x"13"),
  1715 => (x"00",x"00",x"00",x"00"),
  1716 => (x"1a",x"d6",x"00",x"00"),
  1717 => (x"4f",x"42",x"00",x"00"),
  1718 => (x"20",x"20",x"54",x"4f"),
  1719 => (x"4f",x"52",x"20",x"20"),
  1720 => (x"fe",x"1e",x"00",x"4d"),
  1721 => (x"78",x"c0",x"48",x"f0"),
  1722 => (x"09",x"79",x"09",x"cd"),
  1723 => (x"1e",x"1e",x"4f",x"26"),
  1724 => (x"7e",x"bf",x"f0",x"fe"),
  1725 => (x"4f",x"26",x"26",x"48"),
  1726 => (x"48",x"f0",x"fe",x"1e"),
  1727 => (x"4f",x"26",x"78",x"c1"),
  1728 => (x"48",x"f0",x"fe",x"1e"),
  1729 => (x"4f",x"26",x"78",x"c0"),
  1730 => (x"c0",x"4a",x"71",x"1e"),
  1731 => (x"4f",x"26",x"52",x"52"),
  1732 => (x"5c",x"5b",x"5e",x"0e"),
  1733 => (x"86",x"f4",x"0e",x"5d"),
  1734 => (x"6d",x"97",x"4d",x"71"),
  1735 => (x"4c",x"a5",x"c1",x"7e"),
  1736 => (x"c8",x"48",x"6c",x"97"),
  1737 => (x"48",x"6e",x"58",x"a6"),
  1738 => (x"05",x"a8",x"66",x"c4"),
  1739 => (x"48",x"ff",x"87",x"c5"),
  1740 => (x"ff",x"87",x"e6",x"c0"),
  1741 => (x"a5",x"c2",x"87",x"ca"),
  1742 => (x"4b",x"6c",x"97",x"49"),
  1743 => (x"97",x"4b",x"a3",x"71"),
  1744 => (x"6c",x"97",x"4b",x"6b"),
  1745 => (x"c1",x"48",x"6e",x"7e"),
  1746 => (x"58",x"a6",x"c8",x"80"),
  1747 => (x"a6",x"cc",x"98",x"c7"),
  1748 => (x"7c",x"97",x"70",x"58"),
  1749 => (x"73",x"87",x"e1",x"fe"),
  1750 => (x"26",x"8e",x"f4",x"48"),
  1751 => (x"26",x"4c",x"26",x"4d"),
  1752 => (x"0e",x"4f",x"26",x"4b"),
  1753 => (x"0e",x"5c",x"5b",x"5e"),
  1754 => (x"4c",x"71",x"86",x"f4"),
  1755 => (x"c3",x"4a",x"66",x"d8"),
  1756 => (x"a4",x"c2",x"9a",x"ff"),
  1757 => (x"49",x"6c",x"97",x"4b"),
  1758 => (x"72",x"49",x"a1",x"73"),
  1759 => (x"7e",x"6c",x"97",x"51"),
  1760 => (x"80",x"c1",x"48",x"6e"),
  1761 => (x"c7",x"58",x"a6",x"c8"),
  1762 => (x"58",x"a6",x"cc",x"98"),
  1763 => (x"8e",x"f4",x"54",x"70"),
  1764 => (x"1e",x"87",x"ca",x"ff"),
  1765 => (x"87",x"e8",x"fd",x"1e"),
  1766 => (x"49",x"4a",x"bf",x"e0"),
  1767 => (x"99",x"c0",x"e0",x"c0"),
  1768 => (x"72",x"87",x"cb",x"02"),
  1769 => (x"e6",x"f7",x"c2",x"1e"),
  1770 => (x"87",x"f7",x"fe",x"49"),
  1771 => (x"fd",x"fc",x"86",x"c4"),
  1772 => (x"fd",x"7e",x"70",x"87"),
  1773 => (x"26",x"26",x"87",x"c2"),
  1774 => (x"f7",x"c2",x"1e",x"4f"),
  1775 => (x"c7",x"fd",x"49",x"e6"),
  1776 => (x"d3",x"ee",x"c1",x"87"),
  1777 => (x"87",x"da",x"fc",x"49"),
  1778 => (x"26",x"87",x"f7",x"c3"),
  1779 => (x"5b",x"5e",x"0e",x"4f"),
  1780 => (x"71",x"0e",x"5d",x"5c"),
  1781 => (x"e6",x"f7",x"c2",x"4d"),
  1782 => (x"87",x"f4",x"fc",x"49"),
  1783 => (x"b7",x"c0",x"4b",x"70"),
  1784 => (x"c2",x"c3",x"04",x"ab"),
  1785 => (x"ab",x"f0",x"c3",x"87"),
  1786 => (x"c1",x"87",x"c9",x"05"),
  1787 => (x"c1",x"48",x"f1",x"f2"),
  1788 => (x"87",x"e3",x"c2",x"78"),
  1789 => (x"05",x"ab",x"e0",x"c3"),
  1790 => (x"f2",x"c1",x"87",x"c9"),
  1791 => (x"78",x"c1",x"48",x"f5"),
  1792 => (x"c1",x"87",x"d4",x"c2"),
  1793 => (x"02",x"bf",x"f5",x"f2"),
  1794 => (x"c0",x"c2",x"87",x"c6"),
  1795 => (x"87",x"c2",x"4c",x"a3"),
  1796 => (x"f2",x"c1",x"4c",x"73"),
  1797 => (x"c0",x"02",x"bf",x"f1"),
  1798 => (x"49",x"74",x"87",x"e0"),
  1799 => (x"91",x"29",x"b7",x"c4"),
  1800 => (x"81",x"d1",x"f4",x"c1"),
  1801 => (x"9a",x"cf",x"4a",x"74"),
  1802 => (x"48",x"c1",x"92",x"c2"),
  1803 => (x"4a",x"70",x"30",x"72"),
  1804 => (x"48",x"72",x"ba",x"ff"),
  1805 => (x"79",x"70",x"98",x"69"),
  1806 => (x"49",x"74",x"87",x"db"),
  1807 => (x"91",x"29",x"b7",x"c4"),
  1808 => (x"81",x"d1",x"f4",x"c1"),
  1809 => (x"9a",x"cf",x"4a",x"74"),
  1810 => (x"48",x"c3",x"92",x"c2"),
  1811 => (x"4a",x"70",x"30",x"72"),
  1812 => (x"70",x"b0",x"69",x"48"),
  1813 => (x"05",x"9d",x"75",x"79"),
  1814 => (x"ff",x"87",x"f0",x"c0"),
  1815 => (x"e1",x"c8",x"48",x"d0"),
  1816 => (x"48",x"d4",x"ff",x"78"),
  1817 => (x"f2",x"c1",x"78",x"c5"),
  1818 => (x"c3",x"02",x"bf",x"f5"),
  1819 => (x"78",x"e0",x"c3",x"87"),
  1820 => (x"bf",x"f1",x"f2",x"c1"),
  1821 => (x"ff",x"87",x"c6",x"02"),
  1822 => (x"f0",x"c3",x"48",x"d4"),
  1823 => (x"48",x"d4",x"ff",x"78"),
  1824 => (x"d0",x"ff",x"78",x"73"),
  1825 => (x"78",x"e1",x"c8",x"48"),
  1826 => (x"c1",x"78",x"e0",x"c0"),
  1827 => (x"c0",x"48",x"f5",x"f2"),
  1828 => (x"f1",x"f2",x"c1",x"78"),
  1829 => (x"c2",x"78",x"c0",x"48"),
  1830 => (x"f9",x"49",x"e6",x"f7"),
  1831 => (x"4b",x"70",x"87",x"f2"),
  1832 => (x"03",x"ab",x"b7",x"c0"),
  1833 => (x"c0",x"87",x"fe",x"fc"),
  1834 => (x"26",x"4d",x"26",x"48"),
  1835 => (x"26",x"4b",x"26",x"4c"),
  1836 => (x"00",x"00",x"00",x"4f"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"4a",x"71",x"1e",x"00"),
  1839 => (x"87",x"cd",x"fc",x"49"),
  1840 => (x"c0",x"1e",x"4f",x"26"),
  1841 => (x"c4",x"49",x"72",x"4a"),
  1842 => (x"d1",x"f4",x"c1",x"91"),
  1843 => (x"c1",x"79",x"c0",x"81"),
  1844 => (x"aa",x"b7",x"d0",x"82"),
  1845 => (x"26",x"87",x"ee",x"04"),
  1846 => (x"5b",x"5e",x"0e",x"4f"),
  1847 => (x"71",x"0e",x"5d",x"5c"),
  1848 => (x"87",x"dc",x"f8",x"4d"),
  1849 => (x"b7",x"c4",x"4a",x"75"),
  1850 => (x"f4",x"c1",x"92",x"2a"),
  1851 => (x"4c",x"75",x"82",x"d1"),
  1852 => (x"94",x"c2",x"9c",x"cf"),
  1853 => (x"74",x"4b",x"49",x"6a"),
  1854 => (x"c2",x"9b",x"c3",x"2b"),
  1855 => (x"70",x"30",x"74",x"48"),
  1856 => (x"74",x"bc",x"ff",x"4c"),
  1857 => (x"70",x"98",x"71",x"48"),
  1858 => (x"87",x"ec",x"f7",x"7a"),
  1859 => (x"d8",x"fe",x"48",x"73"),
  1860 => (x"00",x"00",x"00",x"87"),
  1861 => (x"00",x"00",x"00",x"00"),
  1862 => (x"00",x"00",x"00",x"00"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"00",x"00"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"00",x"00",x"00",x"00"),
  1868 => (x"00",x"00",x"00",x"00"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"00",x"00"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"d0",x"ff",x"1e",x"00"),
  1877 => (x"78",x"e1",x"c8",x"48"),
  1878 => (x"d4",x"ff",x"48",x"71"),
  1879 => (x"4f",x"26",x"78",x"08"),
  1880 => (x"48",x"d0",x"ff",x"1e"),
  1881 => (x"71",x"78",x"e1",x"c8"),
  1882 => (x"08",x"d4",x"ff",x"48"),
  1883 => (x"48",x"66",x"c4",x"78"),
  1884 => (x"78",x"08",x"d4",x"ff"),
  1885 => (x"71",x"1e",x"4f",x"26"),
  1886 => (x"49",x"66",x"c4",x"4a"),
  1887 => (x"ff",x"49",x"72",x"1e"),
  1888 => (x"d0",x"ff",x"87",x"de"),
  1889 => (x"78",x"e0",x"c0",x"48"),
  1890 => (x"1e",x"4f",x"26",x"26"),
  1891 => (x"4b",x"71",x"1e",x"73"),
  1892 => (x"1e",x"49",x"66",x"c8"),
  1893 => (x"e0",x"c1",x"4a",x"73"),
  1894 => (x"d9",x"ff",x"49",x"a2"),
  1895 => (x"87",x"c4",x"26",x"87"),
  1896 => (x"4c",x"26",x"4d",x"26"),
  1897 => (x"4f",x"26",x"4b",x"26"),
  1898 => (x"71",x"1e",x"73",x"1e"),
  1899 => (x"b7",x"c2",x"4b",x"4a"),
  1900 => (x"87",x"c8",x"03",x"ab"),
  1901 => (x"c3",x"4a",x"49",x"a3"),
  1902 => (x"87",x"c7",x"9a",x"ff"),
  1903 => (x"4a",x"49",x"a3",x"ce"),
  1904 => (x"c8",x"9a",x"ff",x"c3"),
  1905 => (x"72",x"1e",x"49",x"66"),
  1906 => (x"87",x"ea",x"fe",x"49"),
  1907 => (x"87",x"d4",x"ff",x"26"),
  1908 => (x"4a",x"d4",x"ff",x"1e"),
  1909 => (x"ff",x"7a",x"ff",x"c3"),
  1910 => (x"e1",x"c0",x"48",x"d0"),
  1911 => (x"c2",x"7a",x"de",x"78"),
  1912 => (x"7a",x"bf",x"f0",x"f7"),
  1913 => (x"28",x"c8",x"48",x"49"),
  1914 => (x"48",x"71",x"7a",x"70"),
  1915 => (x"7a",x"70",x"28",x"d0"),
  1916 => (x"28",x"d8",x"48",x"71"),
  1917 => (x"d0",x"ff",x"7a",x"70"),
  1918 => (x"78",x"e0",x"c0",x"48"),
  1919 => (x"ff",x"1e",x"4f",x"26"),
  1920 => (x"c9",x"c8",x"48",x"d0"),
  1921 => (x"ff",x"48",x"71",x"78"),
  1922 => (x"26",x"78",x"08",x"d4"),
  1923 => (x"4a",x"71",x"1e",x"4f"),
  1924 => (x"ff",x"87",x"eb",x"49"),
  1925 => (x"78",x"c8",x"48",x"d0"),
  1926 => (x"73",x"1e",x"4f",x"26"),
  1927 => (x"c2",x"4b",x"71",x"1e"),
  1928 => (x"02",x"bf",x"c0",x"f8"),
  1929 => (x"eb",x"c2",x"87",x"c3"),
  1930 => (x"48",x"d0",x"ff",x"87"),
  1931 => (x"73",x"78",x"c9",x"c8"),
  1932 => (x"b1",x"e0",x"c0",x"49"),
  1933 => (x"71",x"48",x"d4",x"ff"),
  1934 => (x"f4",x"f7",x"c2",x"78"),
  1935 => (x"c8",x"78",x"c0",x"48"),
  1936 => (x"87",x"c5",x"02",x"66"),
  1937 => (x"c2",x"49",x"ff",x"c3"),
  1938 => (x"c2",x"49",x"c0",x"87"),
  1939 => (x"cc",x"59",x"fc",x"f7"),
  1940 => (x"87",x"c6",x"02",x"66"),
  1941 => (x"4a",x"d5",x"d5",x"c5"),
  1942 => (x"ff",x"cf",x"87",x"c4"),
  1943 => (x"f8",x"c2",x"4a",x"ff"),
  1944 => (x"f8",x"c2",x"5a",x"c0"),
  1945 => (x"78",x"c1",x"48",x"c0"),
  1946 => (x"4d",x"26",x"87",x"c4"),
  1947 => (x"4b",x"26",x"4c",x"26"),
  1948 => (x"5e",x"0e",x"4f",x"26"),
  1949 => (x"0e",x"5d",x"5c",x"5b"),
  1950 => (x"f7",x"c2",x"4a",x"71"),
  1951 => (x"72",x"4c",x"bf",x"fc"),
  1952 => (x"87",x"cb",x"02",x"9a"),
  1953 => (x"c1",x"91",x"c8",x"49"),
  1954 => (x"71",x"4b",x"d0",x"f8"),
  1955 => (x"c1",x"87",x"c4",x"83"),
  1956 => (x"c0",x"4b",x"d0",x"fc"),
  1957 => (x"74",x"49",x"13",x"4d"),
  1958 => (x"f8",x"f7",x"c2",x"99"),
  1959 => (x"d4",x"ff",x"b9",x"bf"),
  1960 => (x"c1",x"78",x"71",x"48"),
  1961 => (x"c8",x"85",x"2c",x"b7"),
  1962 => (x"e8",x"04",x"ad",x"b7"),
  1963 => (x"f4",x"f7",x"c2",x"87"),
  1964 => (x"80",x"c8",x"48",x"bf"),
  1965 => (x"58",x"f8",x"f7",x"c2"),
  1966 => (x"1e",x"87",x"ef",x"fe"),
  1967 => (x"4b",x"71",x"1e",x"73"),
  1968 => (x"02",x"9a",x"4a",x"13"),
  1969 => (x"49",x"72",x"87",x"cb"),
  1970 => (x"13",x"87",x"e7",x"fe"),
  1971 => (x"f5",x"05",x"9a",x"4a"),
  1972 => (x"87",x"da",x"fe",x"87"),
  1973 => (x"f4",x"f7",x"c2",x"1e"),
  1974 => (x"f7",x"c2",x"49",x"bf"),
  1975 => (x"a1",x"c1",x"48",x"f4"),
  1976 => (x"b7",x"c0",x"c4",x"78"),
  1977 => (x"87",x"db",x"03",x"a9"),
  1978 => (x"c2",x"48",x"d4",x"ff"),
  1979 => (x"78",x"bf",x"f8",x"f7"),
  1980 => (x"bf",x"f4",x"f7",x"c2"),
  1981 => (x"f4",x"f7",x"c2",x"49"),
  1982 => (x"78",x"a1",x"c1",x"48"),
  1983 => (x"a9",x"b7",x"c0",x"c4"),
  1984 => (x"ff",x"87",x"e5",x"04"),
  1985 => (x"78",x"c8",x"48",x"d0"),
  1986 => (x"48",x"c0",x"f8",x"c2"),
  1987 => (x"4f",x"26",x"78",x"c0"),
  1988 => (x"00",x"00",x"00",x"00"),
  1989 => (x"00",x"00",x"00",x"00"),
  1990 => (x"5f",x"00",x"00",x"00"),
  1991 => (x"00",x"00",x"00",x"5f"),
  1992 => (x"00",x"03",x"03",x"00"),
  1993 => (x"00",x"00",x"03",x"03"),
  1994 => (x"14",x"7f",x"7f",x"14"),
  1995 => (x"00",x"14",x"7f",x"7f"),
  1996 => (x"6b",x"2e",x"24",x"00"),
  1997 => (x"00",x"12",x"3a",x"6b"),
  1998 => (x"18",x"36",x"6a",x"4c"),
  1999 => (x"00",x"32",x"56",x"6c"),
  2000 => (x"59",x"4f",x"7e",x"30"),
  2001 => (x"40",x"68",x"3a",x"77"),
  2002 => (x"07",x"04",x"00",x"00"),
  2003 => (x"00",x"00",x"00",x"03"),
  2004 => (x"3e",x"1c",x"00",x"00"),
  2005 => (x"00",x"00",x"41",x"63"),
  2006 => (x"63",x"41",x"00",x"00"),
  2007 => (x"00",x"00",x"1c",x"3e"),
  2008 => (x"1c",x"3e",x"2a",x"08"),
  2009 => (x"08",x"2a",x"3e",x"1c"),
  2010 => (x"3e",x"08",x"08",x"00"),
  2011 => (x"00",x"08",x"08",x"3e"),
  2012 => (x"e0",x"80",x"00",x"00"),
  2013 => (x"00",x"00",x"00",x"60"),
  2014 => (x"08",x"08",x"08",x"00"),
  2015 => (x"00",x"08",x"08",x"08"),
  2016 => (x"60",x"00",x"00",x"00"),
  2017 => (x"00",x"00",x"00",x"60"),
  2018 => (x"18",x"30",x"60",x"40"),
  2019 => (x"01",x"03",x"06",x"0c"),
  2020 => (x"59",x"7f",x"3e",x"00"),
  2021 => (x"00",x"3e",x"7f",x"4d"),
  2022 => (x"7f",x"06",x"04",x"00"),
  2023 => (x"00",x"00",x"00",x"7f"),
  2024 => (x"71",x"63",x"42",x"00"),
  2025 => (x"00",x"46",x"4f",x"59"),
  2026 => (x"49",x"63",x"22",x"00"),
  2027 => (x"00",x"36",x"7f",x"49"),
  2028 => (x"13",x"16",x"1c",x"18"),
  2029 => (x"00",x"10",x"7f",x"7f"),
  2030 => (x"45",x"67",x"27",x"00"),
  2031 => (x"00",x"39",x"7d",x"45"),
  2032 => (x"4b",x"7e",x"3c",x"00"),
  2033 => (x"00",x"30",x"79",x"49"),
  2034 => (x"71",x"01",x"01",x"00"),
  2035 => (x"00",x"07",x"0f",x"79"),
  2036 => (x"49",x"7f",x"36",x"00"),
  2037 => (x"00",x"36",x"7f",x"49"),
  2038 => (x"49",x"4f",x"06",x"00"),
  2039 => (x"00",x"1e",x"3f",x"69"),
  2040 => (x"66",x"00",x"00",x"00"),
  2041 => (x"00",x"00",x"00",x"66"),
  2042 => (x"e6",x"80",x"00",x"00"),
  2043 => (x"00",x"00",x"00",x"66"),
  2044 => (x"14",x"08",x"08",x"00"),
  2045 => (x"00",x"22",x"22",x"14"),
  2046 => (x"14",x"14",x"14",x"00"),
  2047 => (x"00",x"14",x"14",x"14"),
  2048 => (x"14",x"22",x"22",x"00"),
  2049 => (x"00",x"08",x"08",x"14"),
  2050 => (x"51",x"03",x"02",x"00"),
  2051 => (x"00",x"06",x"0f",x"59"),
  2052 => (x"5d",x"41",x"7f",x"3e"),
  2053 => (x"00",x"1e",x"1f",x"55"),
  2054 => (x"09",x"7f",x"7e",x"00"),
  2055 => (x"00",x"7e",x"7f",x"09"),
  2056 => (x"49",x"7f",x"7f",x"00"),
  2057 => (x"00",x"36",x"7f",x"49"),
  2058 => (x"63",x"3e",x"1c",x"00"),
  2059 => (x"00",x"41",x"41",x"41"),
  2060 => (x"41",x"7f",x"7f",x"00"),
  2061 => (x"00",x"1c",x"3e",x"63"),
  2062 => (x"49",x"7f",x"7f",x"00"),
  2063 => (x"00",x"41",x"41",x"49"),
  2064 => (x"09",x"7f",x"7f",x"00"),
  2065 => (x"00",x"01",x"01",x"09"),
  2066 => (x"41",x"7f",x"3e",x"00"),
  2067 => (x"00",x"7a",x"7b",x"49"),
  2068 => (x"08",x"7f",x"7f",x"00"),
  2069 => (x"00",x"7f",x"7f",x"08"),
  2070 => (x"7f",x"41",x"00",x"00"),
  2071 => (x"00",x"00",x"41",x"7f"),
  2072 => (x"40",x"60",x"20",x"00"),
  2073 => (x"00",x"3f",x"7f",x"40"),
  2074 => (x"1c",x"08",x"7f",x"7f"),
  2075 => (x"00",x"41",x"63",x"36"),
  2076 => (x"40",x"7f",x"7f",x"00"),
  2077 => (x"00",x"40",x"40",x"40"),
  2078 => (x"0c",x"06",x"7f",x"7f"),
  2079 => (x"00",x"7f",x"7f",x"06"),
  2080 => (x"0c",x"06",x"7f",x"7f"),
  2081 => (x"00",x"7f",x"7f",x"18"),
  2082 => (x"41",x"7f",x"3e",x"00"),
  2083 => (x"00",x"3e",x"7f",x"41"),
  2084 => (x"09",x"7f",x"7f",x"00"),
  2085 => (x"00",x"06",x"0f",x"09"),
  2086 => (x"61",x"41",x"7f",x"3e"),
  2087 => (x"00",x"40",x"7e",x"7f"),
  2088 => (x"09",x"7f",x"7f",x"00"),
  2089 => (x"00",x"66",x"7f",x"19"),
  2090 => (x"4d",x"6f",x"26",x"00"),
  2091 => (x"00",x"32",x"7b",x"59"),
  2092 => (x"7f",x"01",x"01",x"00"),
  2093 => (x"00",x"01",x"01",x"7f"),
  2094 => (x"40",x"7f",x"3f",x"00"),
  2095 => (x"00",x"3f",x"7f",x"40"),
  2096 => (x"70",x"3f",x"0f",x"00"),
  2097 => (x"00",x"0f",x"3f",x"70"),
  2098 => (x"18",x"30",x"7f",x"7f"),
  2099 => (x"00",x"7f",x"7f",x"30"),
  2100 => (x"1c",x"36",x"63",x"41"),
  2101 => (x"41",x"63",x"36",x"1c"),
  2102 => (x"7c",x"06",x"03",x"01"),
  2103 => (x"01",x"03",x"06",x"7c"),
  2104 => (x"4d",x"59",x"71",x"61"),
  2105 => (x"00",x"41",x"43",x"47"),
  2106 => (x"7f",x"7f",x"00",x"00"),
  2107 => (x"00",x"00",x"41",x"41"),
  2108 => (x"0c",x"06",x"03",x"01"),
  2109 => (x"40",x"60",x"30",x"18"),
  2110 => (x"41",x"41",x"00",x"00"),
  2111 => (x"00",x"00",x"7f",x"7f"),
  2112 => (x"03",x"06",x"0c",x"08"),
  2113 => (x"00",x"08",x"0c",x"06"),
  2114 => (x"80",x"80",x"80",x"80"),
  2115 => (x"00",x"80",x"80",x"80"),
  2116 => (x"03",x"00",x"00",x"00"),
  2117 => (x"00",x"00",x"04",x"07"),
  2118 => (x"54",x"74",x"20",x"00"),
  2119 => (x"00",x"78",x"7c",x"54"),
  2120 => (x"44",x"7f",x"7f",x"00"),
  2121 => (x"00",x"38",x"7c",x"44"),
  2122 => (x"44",x"7c",x"38",x"00"),
  2123 => (x"00",x"00",x"44",x"44"),
  2124 => (x"44",x"7c",x"38",x"00"),
  2125 => (x"00",x"7f",x"7f",x"44"),
  2126 => (x"54",x"7c",x"38",x"00"),
  2127 => (x"00",x"18",x"5c",x"54"),
  2128 => (x"7f",x"7e",x"04",x"00"),
  2129 => (x"00",x"00",x"05",x"05"),
  2130 => (x"a4",x"bc",x"18",x"00"),
  2131 => (x"00",x"7c",x"fc",x"a4"),
  2132 => (x"04",x"7f",x"7f",x"00"),
  2133 => (x"00",x"78",x"7c",x"04"),
  2134 => (x"3d",x"00",x"00",x"00"),
  2135 => (x"00",x"00",x"40",x"7d"),
  2136 => (x"80",x"80",x"80",x"00"),
  2137 => (x"00",x"00",x"7d",x"fd"),
  2138 => (x"10",x"7f",x"7f",x"00"),
  2139 => (x"00",x"44",x"6c",x"38"),
  2140 => (x"3f",x"00",x"00",x"00"),
  2141 => (x"00",x"00",x"40",x"7f"),
  2142 => (x"18",x"0c",x"7c",x"7c"),
  2143 => (x"00",x"78",x"7c",x"0c"),
  2144 => (x"04",x"7c",x"7c",x"00"),
  2145 => (x"00",x"78",x"7c",x"04"),
  2146 => (x"44",x"7c",x"38",x"00"),
  2147 => (x"00",x"38",x"7c",x"44"),
  2148 => (x"24",x"fc",x"fc",x"00"),
  2149 => (x"00",x"18",x"3c",x"24"),
  2150 => (x"24",x"3c",x"18",x"00"),
  2151 => (x"00",x"fc",x"fc",x"24"),
  2152 => (x"04",x"7c",x"7c",x"00"),
  2153 => (x"00",x"08",x"0c",x"04"),
  2154 => (x"54",x"5c",x"48",x"00"),
  2155 => (x"00",x"20",x"74",x"54"),
  2156 => (x"7f",x"3f",x"04",x"00"),
  2157 => (x"00",x"00",x"44",x"44"),
  2158 => (x"40",x"7c",x"3c",x"00"),
  2159 => (x"00",x"7c",x"7c",x"40"),
  2160 => (x"60",x"3c",x"1c",x"00"),
  2161 => (x"00",x"1c",x"3c",x"60"),
  2162 => (x"30",x"60",x"7c",x"3c"),
  2163 => (x"00",x"3c",x"7c",x"60"),
  2164 => (x"10",x"38",x"6c",x"44"),
  2165 => (x"00",x"44",x"6c",x"38"),
  2166 => (x"e0",x"bc",x"1c",x"00"),
  2167 => (x"00",x"1c",x"3c",x"60"),
  2168 => (x"74",x"64",x"44",x"00"),
  2169 => (x"00",x"44",x"4c",x"5c"),
  2170 => (x"3e",x"08",x"08",x"00"),
  2171 => (x"00",x"41",x"41",x"77"),
  2172 => (x"7f",x"00",x"00",x"00"),
  2173 => (x"00",x"00",x"00",x"7f"),
  2174 => (x"77",x"41",x"41",x"00"),
  2175 => (x"00",x"08",x"08",x"3e"),
  2176 => (x"03",x"01",x"01",x"02"),
  2177 => (x"00",x"01",x"02",x"02"),
  2178 => (x"7f",x"7f",x"7f",x"7f"),
  2179 => (x"00",x"7f",x"7f",x"7f"),
  2180 => (x"1c",x"1c",x"08",x"08"),
  2181 => (x"7f",x"7f",x"3e",x"3e"),
  2182 => (x"3e",x"3e",x"7f",x"7f"),
  2183 => (x"08",x"08",x"1c",x"1c"),
  2184 => (x"7c",x"18",x"10",x"00"),
  2185 => (x"00",x"10",x"18",x"7c"),
  2186 => (x"7c",x"30",x"10",x"00"),
  2187 => (x"00",x"10",x"30",x"7c"),
  2188 => (x"60",x"60",x"30",x"10"),
  2189 => (x"00",x"06",x"1e",x"78"),
  2190 => (x"18",x"3c",x"66",x"42"),
  2191 => (x"00",x"42",x"66",x"3c"),
  2192 => (x"c2",x"6a",x"38",x"78"),
  2193 => (x"00",x"38",x"6c",x"c6"),
  2194 => (x"60",x"00",x"00",x"60"),
  2195 => (x"00",x"60",x"00",x"00"),
  2196 => (x"5c",x"5b",x"5e",x"0e"),
  2197 => (x"71",x"1e",x"0e",x"5d"),
  2198 => (x"d1",x"f8",x"c2",x"4c"),
  2199 => (x"4b",x"c0",x"4d",x"bf"),
  2200 => (x"ab",x"74",x"1e",x"c0"),
  2201 => (x"c4",x"87",x"c7",x"02"),
  2202 => (x"78",x"c0",x"48",x"a6"),
  2203 => (x"a6",x"c4",x"87",x"c5"),
  2204 => (x"c4",x"78",x"c1",x"48"),
  2205 => (x"49",x"73",x"1e",x"66"),
  2206 => (x"c8",x"87",x"df",x"ee"),
  2207 => (x"49",x"e0",x"c0",x"86"),
  2208 => (x"c4",x"87",x"ef",x"ef"),
  2209 => (x"49",x"6a",x"4a",x"a5"),
  2210 => (x"f1",x"87",x"f0",x"f0"),
  2211 => (x"85",x"cb",x"87",x"c6"),
  2212 => (x"b7",x"c8",x"83",x"c1"),
  2213 => (x"c7",x"ff",x"04",x"ab"),
  2214 => (x"4d",x"26",x"26",x"87"),
  2215 => (x"4b",x"26",x"4c",x"26"),
  2216 => (x"71",x"1e",x"4f",x"26"),
  2217 => (x"d5",x"f8",x"c2",x"4a"),
  2218 => (x"d5",x"f8",x"c2",x"5a"),
  2219 => (x"49",x"78",x"c7",x"48"),
  2220 => (x"26",x"87",x"dd",x"fe"),
  2221 => (x"1e",x"73",x"1e",x"4f"),
  2222 => (x"b7",x"c0",x"4a",x"71"),
  2223 => (x"87",x"d3",x"03",x"aa"),
  2224 => (x"bf",x"f6",x"db",x"c2"),
  2225 => (x"c1",x"87",x"c4",x"05"),
  2226 => (x"c0",x"87",x"c2",x"4b"),
  2227 => (x"fa",x"db",x"c2",x"4b"),
  2228 => (x"c2",x"87",x"c4",x"5b"),
  2229 => (x"c2",x"5a",x"fa",x"db"),
  2230 => (x"4a",x"bf",x"f6",x"db"),
  2231 => (x"c0",x"c1",x"9a",x"c1"),
  2232 => (x"e8",x"ec",x"49",x"a2"),
  2233 => (x"de",x"db",x"c2",x"87"),
  2234 => (x"db",x"c2",x"49",x"bf"),
  2235 => (x"fc",x"b1",x"bf",x"f6"),
  2236 => (x"fe",x"78",x"71",x"48"),
  2237 => (x"71",x"1e",x"87",x"e8"),
  2238 => (x"1e",x"66",x"c4",x"4a"),
  2239 => (x"e7",x"ea",x"49",x"72"),
  2240 => (x"4f",x"26",x"26",x"87"),
  2241 => (x"ff",x"4a",x"71",x"1e"),
  2242 => (x"ff",x"c3",x"48",x"d4"),
  2243 => (x"48",x"d0",x"ff",x"78"),
  2244 => (x"ff",x"78",x"e1",x"c0"),
  2245 => (x"78",x"c1",x"48",x"d4"),
  2246 => (x"31",x"c4",x"49",x"72"),
  2247 => (x"d0",x"ff",x"78",x"71"),
  2248 => (x"78",x"e0",x"c0",x"48"),
  2249 => (x"c2",x"1e",x"4f",x"26"),
  2250 => (x"49",x"bf",x"f6",x"db"),
  2251 => (x"c2",x"87",x"ca",x"e6"),
  2252 => (x"e8",x"48",x"c9",x"f8"),
  2253 => (x"f8",x"c2",x"78",x"bf"),
  2254 => (x"bf",x"ec",x"48",x"c5"),
  2255 => (x"c9",x"f8",x"c2",x"78"),
  2256 => (x"c3",x"49",x"4a",x"bf"),
  2257 => (x"b7",x"c8",x"99",x"ff"),
  2258 => (x"71",x"48",x"72",x"2a"),
  2259 => (x"d1",x"f8",x"c2",x"b0"),
  2260 => (x"0e",x"4f",x"26",x"58"),
  2261 => (x"5d",x"5c",x"5b",x"5e"),
  2262 => (x"ff",x"4b",x"71",x"0e"),
  2263 => (x"f8",x"c2",x"87",x"c8"),
  2264 => (x"50",x"c0",x"48",x"c4"),
  2265 => (x"f0",x"e5",x"49",x"73"),
  2266 => (x"4c",x"49",x"70",x"87"),
  2267 => (x"ee",x"cb",x"9c",x"c2"),
  2268 => (x"87",x"ca",x"ce",x"49"),
  2269 => (x"c2",x"4d",x"49",x"70"),
  2270 => (x"bf",x"97",x"c4",x"f8"),
  2271 => (x"87",x"e2",x"c1",x"05"),
  2272 => (x"c2",x"49",x"66",x"d0"),
  2273 => (x"99",x"bf",x"cd",x"f8"),
  2274 => (x"d4",x"87",x"d6",x"05"),
  2275 => (x"f8",x"c2",x"49",x"66"),
  2276 => (x"05",x"99",x"bf",x"c5"),
  2277 => (x"49",x"73",x"87",x"cb"),
  2278 => (x"70",x"87",x"fe",x"e4"),
  2279 => (x"c1",x"c1",x"02",x"98"),
  2280 => (x"fe",x"4c",x"c1",x"87"),
  2281 => (x"49",x"75",x"87",x"c0"),
  2282 => (x"70",x"87",x"df",x"cd"),
  2283 => (x"87",x"c6",x"02",x"98"),
  2284 => (x"48",x"c4",x"f8",x"c2"),
  2285 => (x"f8",x"c2",x"50",x"c1"),
  2286 => (x"05",x"bf",x"97",x"c4"),
  2287 => (x"c2",x"87",x"e3",x"c0"),
  2288 => (x"49",x"bf",x"cd",x"f8"),
  2289 => (x"05",x"99",x"66",x"d0"),
  2290 => (x"c2",x"87",x"d6",x"ff"),
  2291 => (x"49",x"bf",x"c5",x"f8"),
  2292 => (x"05",x"99",x"66",x"d4"),
  2293 => (x"73",x"87",x"ca",x"ff"),
  2294 => (x"87",x"fd",x"e3",x"49"),
  2295 => (x"fe",x"05",x"98",x"70"),
  2296 => (x"48",x"74",x"87",x"ff"),
  2297 => (x"0e",x"87",x"f3",x"fa"),
  2298 => (x"5d",x"5c",x"5b",x"5e"),
  2299 => (x"c0",x"86",x"f4",x"0e"),
  2300 => (x"bf",x"ec",x"4c",x"4d"),
  2301 => (x"48",x"a6",x"c4",x"7e"),
  2302 => (x"bf",x"d1",x"f8",x"c2"),
  2303 => (x"1e",x"1e",x"c0",x"78"),
  2304 => (x"fd",x"49",x"f7",x"c1"),
  2305 => (x"86",x"c8",x"87",x"cd"),
  2306 => (x"c0",x"02",x"98",x"70"),
  2307 => (x"db",x"c2",x"87",x"f3"),
  2308 => (x"c4",x"05",x"bf",x"de"),
  2309 => (x"c2",x"7e",x"c1",x"87"),
  2310 => (x"c2",x"7e",x"c0",x"87"),
  2311 => (x"6e",x"48",x"de",x"db"),
  2312 => (x"1e",x"fc",x"ca",x"78"),
  2313 => (x"c9",x"02",x"66",x"c4"),
  2314 => (x"48",x"a6",x"c4",x"87"),
  2315 => (x"78",x"f1",x"d9",x"c2"),
  2316 => (x"a6",x"c4",x"87",x"c7"),
  2317 => (x"fc",x"d9",x"c2",x"48"),
  2318 => (x"49",x"66",x"c4",x"78"),
  2319 => (x"c4",x"87",x"c9",x"c9"),
  2320 => (x"c0",x"1e",x"c1",x"86"),
  2321 => (x"fc",x"49",x"c7",x"1e"),
  2322 => (x"86",x"c8",x"87",x"c9"),
  2323 => (x"cd",x"02",x"98",x"70"),
  2324 => (x"f9",x"49",x"ff",x"87"),
  2325 => (x"da",x"c1",x"87",x"df"),
  2326 => (x"87",x"fd",x"e1",x"49"),
  2327 => (x"f8",x"c2",x"4d",x"c1"),
  2328 => (x"02",x"bf",x"97",x"c4"),
  2329 => (x"db",x"c2",x"87",x"cf"),
  2330 => (x"c1",x"49",x"bf",x"da"),
  2331 => (x"de",x"db",x"c2",x"b9"),
  2332 => (x"cf",x"fa",x"71",x"59"),
  2333 => (x"c9",x"f8",x"c2",x"87"),
  2334 => (x"db",x"c2",x"4b",x"bf"),
  2335 => (x"c1",x"05",x"bf",x"f6"),
  2336 => (x"db",x"c2",x"87",x"e1"),
  2337 => (x"c0",x"02",x"bf",x"de"),
  2338 => (x"a6",x"c4",x"87",x"f0"),
  2339 => (x"c0",x"c0",x"c8",x"48"),
  2340 => (x"e2",x"db",x"c2",x"78"),
  2341 => (x"bf",x"97",x"6e",x"7e"),
  2342 => (x"c1",x"48",x"6e",x"49"),
  2343 => (x"71",x"7e",x"70",x"80"),
  2344 => (x"70",x"87",x"f6",x"e0"),
  2345 => (x"87",x"c3",x"02",x"98"),
  2346 => (x"c4",x"b3",x"66",x"c4"),
  2347 => (x"b7",x"c1",x"48",x"66"),
  2348 => (x"58",x"a6",x"c8",x"28"),
  2349 => (x"ff",x"05",x"98",x"70"),
  2350 => (x"fd",x"c3",x"87",x"db"),
  2351 => (x"87",x"d9",x"e0",x"49"),
  2352 => (x"e0",x"49",x"fa",x"c3"),
  2353 => (x"49",x"73",x"87",x"d3"),
  2354 => (x"71",x"99",x"ff",x"c3"),
  2355 => (x"f8",x"49",x"c0",x"1e"),
  2356 => (x"49",x"73",x"87",x"e4"),
  2357 => (x"71",x"29",x"b7",x"c8"),
  2358 => (x"f8",x"49",x"c1",x"1e"),
  2359 => (x"86",x"c8",x"87",x"d8"),
  2360 => (x"c2",x"87",x"c9",x"c6"),
  2361 => (x"4b",x"bf",x"cd",x"f8"),
  2362 => (x"87",x"df",x"02",x"9b"),
  2363 => (x"bf",x"f2",x"db",x"c2"),
  2364 => (x"87",x"d6",x"c8",x"49"),
  2365 => (x"c0",x"05",x"98",x"70"),
  2366 => (x"4b",x"c0",x"87",x"c4"),
  2367 => (x"e0",x"c2",x"87",x"d3"),
  2368 => (x"87",x"fa",x"c7",x"49"),
  2369 => (x"58",x"f6",x"db",x"c2"),
  2370 => (x"c2",x"87",x"c6",x"c0"),
  2371 => (x"c0",x"48",x"f2",x"db"),
  2372 => (x"c2",x"49",x"73",x"78"),
  2373 => (x"cf",x"c0",x"05",x"99"),
  2374 => (x"49",x"eb",x"c3",x"87"),
  2375 => (x"87",x"f9",x"de",x"ff"),
  2376 => (x"99",x"c2",x"49",x"70"),
  2377 => (x"87",x"c2",x"c0",x"02"),
  2378 => (x"49",x"73",x"4c",x"fb"),
  2379 => (x"c0",x"05",x"99",x"c1"),
  2380 => (x"f4",x"c3",x"87",x"cf"),
  2381 => (x"e0",x"de",x"ff",x"49"),
  2382 => (x"c2",x"49",x"70",x"87"),
  2383 => (x"c2",x"c0",x"02",x"99"),
  2384 => (x"73",x"4c",x"fa",x"87"),
  2385 => (x"05",x"99",x"c8",x"49"),
  2386 => (x"c3",x"87",x"cf",x"c0"),
  2387 => (x"de",x"ff",x"49",x"f5"),
  2388 => (x"49",x"70",x"87",x"c7"),
  2389 => (x"c0",x"02",x"99",x"c2"),
  2390 => (x"f8",x"c2",x"87",x"d6"),
  2391 => (x"c0",x"02",x"bf",x"d5"),
  2392 => (x"c1",x"48",x"87",x"ca"),
  2393 => (x"d9",x"f8",x"c2",x"88"),
  2394 => (x"87",x"c2",x"c0",x"58"),
  2395 => (x"4d",x"c1",x"4c",x"ff"),
  2396 => (x"99",x"c4",x"49",x"73"),
  2397 => (x"87",x"cf",x"c0",x"05"),
  2398 => (x"ff",x"49",x"f2",x"c3"),
  2399 => (x"70",x"87",x"da",x"dd"),
  2400 => (x"02",x"99",x"c2",x"49"),
  2401 => (x"c2",x"87",x"dc",x"c0"),
  2402 => (x"7e",x"bf",x"d5",x"f8"),
  2403 => (x"a8",x"b7",x"c7",x"48"),
  2404 => (x"87",x"cb",x"c0",x"03"),
  2405 => (x"80",x"c1",x"48",x"6e"),
  2406 => (x"58",x"d9",x"f8",x"c2"),
  2407 => (x"fe",x"87",x"c2",x"c0"),
  2408 => (x"c3",x"4d",x"c1",x"4c"),
  2409 => (x"dc",x"ff",x"49",x"fd"),
  2410 => (x"49",x"70",x"87",x"ef"),
  2411 => (x"c0",x"02",x"99",x"c2"),
  2412 => (x"f8",x"c2",x"87",x"d5"),
  2413 => (x"c0",x"02",x"bf",x"d5"),
  2414 => (x"f8",x"c2",x"87",x"c9"),
  2415 => (x"78",x"c0",x"48",x"d5"),
  2416 => (x"fd",x"87",x"c2",x"c0"),
  2417 => (x"c3",x"4d",x"c1",x"4c"),
  2418 => (x"dc",x"ff",x"49",x"fa"),
  2419 => (x"49",x"70",x"87",x"cb"),
  2420 => (x"c0",x"02",x"99",x"c2"),
  2421 => (x"f8",x"c2",x"87",x"d9"),
  2422 => (x"c7",x"48",x"bf",x"d5"),
  2423 => (x"c0",x"03",x"a8",x"b7"),
  2424 => (x"f8",x"c2",x"87",x"c9"),
  2425 => (x"78",x"c7",x"48",x"d5"),
  2426 => (x"fc",x"87",x"c2",x"c0"),
  2427 => (x"c0",x"4d",x"c1",x"4c"),
  2428 => (x"c0",x"03",x"ac",x"b7"),
  2429 => (x"66",x"c4",x"87",x"d0"),
  2430 => (x"82",x"d8",x"c1",x"4a"),
  2431 => (x"c5",x"c0",x"02",x"6a"),
  2432 => (x"49",x"74",x"4b",x"87"),
  2433 => (x"1e",x"c0",x"0f",x"73"),
  2434 => (x"c1",x"1e",x"f0",x"c3"),
  2435 => (x"c2",x"f5",x"49",x"da"),
  2436 => (x"70",x"86",x"c8",x"87"),
  2437 => (x"e0",x"c0",x"02",x"98"),
  2438 => (x"48",x"a6",x"c8",x"87"),
  2439 => (x"bf",x"d5",x"f8",x"c2"),
  2440 => (x"49",x"66",x"c8",x"78"),
  2441 => (x"66",x"c4",x"91",x"cb"),
  2442 => (x"70",x"80",x"71",x"48"),
  2443 => (x"02",x"bf",x"6e",x"7e"),
  2444 => (x"4b",x"87",x"c6",x"c0"),
  2445 => (x"73",x"49",x"66",x"c8"),
  2446 => (x"02",x"9d",x"75",x"0f"),
  2447 => (x"c2",x"87",x"c8",x"c0"),
  2448 => (x"49",x"bf",x"d5",x"f8"),
  2449 => (x"c2",x"87",x"c9",x"f0"),
  2450 => (x"02",x"bf",x"fa",x"db"),
  2451 => (x"49",x"87",x"dd",x"c0"),
  2452 => (x"70",x"87",x"f7",x"c2"),
  2453 => (x"d3",x"c0",x"02",x"98"),
  2454 => (x"d5",x"f8",x"c2",x"87"),
  2455 => (x"ef",x"ef",x"49",x"bf"),
  2456 => (x"f1",x"49",x"c0",x"87"),
  2457 => (x"db",x"c2",x"87",x"cf"),
  2458 => (x"78",x"c0",x"48",x"fa"),
  2459 => (x"e9",x"f0",x"8e",x"f4"),
  2460 => (x"79",x"6f",x"4a",x"87"),
  2461 => (x"73",x"79",x"65",x"6b"),
  2462 => (x"00",x"6e",x"6f",x"20"),
  2463 => (x"6b",x"79",x"6f",x"4a"),
  2464 => (x"20",x"73",x"79",x"65"),
  2465 => (x"00",x"66",x"66",x"6f"),
  2466 => (x"5c",x"5b",x"5e",x"0e"),
  2467 => (x"71",x"1e",x"0e",x"5d"),
  2468 => (x"d1",x"f8",x"c2",x"4c"),
  2469 => (x"cd",x"c1",x"49",x"bf"),
  2470 => (x"d1",x"c1",x"4d",x"a1"),
  2471 => (x"74",x"7e",x"69",x"81"),
  2472 => (x"87",x"cf",x"02",x"9c"),
  2473 => (x"74",x"4b",x"a5",x"c4"),
  2474 => (x"d1",x"f8",x"c2",x"7b"),
  2475 => (x"f1",x"ef",x"49",x"bf"),
  2476 => (x"74",x"7b",x"6e",x"87"),
  2477 => (x"87",x"c4",x"05",x"9c"),
  2478 => (x"87",x"c2",x"4b",x"c0"),
  2479 => (x"49",x"73",x"4b",x"c1"),
  2480 => (x"d4",x"87",x"f2",x"ef"),
  2481 => (x"87",x"c8",x"02",x"66"),
  2482 => (x"87",x"f2",x"c0",x"49"),
  2483 => (x"87",x"c2",x"4a",x"70"),
  2484 => (x"db",x"c2",x"4a",x"c0"),
  2485 => (x"ef",x"26",x"5a",x"fe"),
  2486 => (x"00",x"00",x"87",x"c0"),
  2487 => (x"00",x"00",x"00",x"00"),
  2488 => (x"12",x"58",x"00",x"00"),
  2489 => (x"1b",x"1d",x"14",x"11"),
  2490 => (x"59",x"5a",x"23",x"1c"),
  2491 => (x"f2",x"f5",x"94",x"91"),
  2492 => (x"00",x"00",x"f4",x"eb"),
  2493 => (x"00",x"00",x"00",x"00"),
  2494 => (x"00",x"00",x"00",x"00"),
  2495 => (x"71",x"1e",x"00",x"00"),
  2496 => (x"bf",x"c8",x"ff",x"4a"),
  2497 => (x"48",x"a1",x"72",x"49"),
  2498 => (x"ff",x"1e",x"4f",x"26"),
  2499 => (x"fe",x"89",x"bf",x"c8"),
  2500 => (x"c0",x"c0",x"c0",x"c0"),
  2501 => (x"c4",x"01",x"a9",x"c0"),
  2502 => (x"c2",x"4a",x"c0",x"87"),
  2503 => (x"72",x"4a",x"c1",x"87"),
  2504 => (x"0e",x"4f",x"26",x"48"),
  2505 => (x"5d",x"5c",x"5b",x"5e"),
  2506 => (x"ff",x"4b",x"71",x"0e"),
  2507 => (x"66",x"d0",x"4c",x"d4"),
  2508 => (x"d6",x"78",x"c0",x"48"),
  2509 => (x"d8",x"d8",x"ff",x"49"),
  2510 => (x"7c",x"ff",x"c3",x"87"),
  2511 => (x"ff",x"c3",x"49",x"6c"),
  2512 => (x"49",x"4d",x"71",x"99"),
  2513 => (x"c1",x"99",x"f0",x"c3"),
  2514 => (x"cb",x"05",x"a9",x"e0"),
  2515 => (x"7c",x"ff",x"c3",x"87"),
  2516 => (x"98",x"c3",x"48",x"6c"),
  2517 => (x"78",x"08",x"66",x"d0"),
  2518 => (x"6c",x"7c",x"ff",x"c3"),
  2519 => (x"31",x"c8",x"49",x"4a"),
  2520 => (x"6c",x"7c",x"ff",x"c3"),
  2521 => (x"72",x"b2",x"71",x"4a"),
  2522 => (x"c3",x"31",x"c8",x"49"),
  2523 => (x"4a",x"6c",x"7c",x"ff"),
  2524 => (x"49",x"72",x"b2",x"71"),
  2525 => (x"ff",x"c3",x"31",x"c8"),
  2526 => (x"71",x"4a",x"6c",x"7c"),
  2527 => (x"48",x"d0",x"ff",x"b2"),
  2528 => (x"73",x"78",x"e0",x"c0"),
  2529 => (x"87",x"c2",x"02",x"9b"),
  2530 => (x"48",x"75",x"7b",x"72"),
  2531 => (x"4c",x"26",x"4d",x"26"),
  2532 => (x"4f",x"26",x"4b",x"26"),
  2533 => (x"0e",x"4f",x"26",x"1e"),
  2534 => (x"0e",x"5c",x"5b",x"5e"),
  2535 => (x"1e",x"76",x"86",x"f8"),
  2536 => (x"fd",x"49",x"a6",x"c8"),
  2537 => (x"86",x"c4",x"87",x"fd"),
  2538 => (x"48",x"6e",x"4b",x"70"),
  2539 => (x"c2",x"03",x"a8",x"c2"),
  2540 => (x"4a",x"73",x"87",x"f0"),
  2541 => (x"c1",x"9a",x"f0",x"c3"),
  2542 => (x"c7",x"02",x"aa",x"d0"),
  2543 => (x"aa",x"e0",x"c1",x"87"),
  2544 => (x"87",x"de",x"c2",x"05"),
  2545 => (x"99",x"c8",x"49",x"73"),
  2546 => (x"ff",x"87",x"c3",x"02"),
  2547 => (x"4c",x"73",x"87",x"c6"),
  2548 => (x"ac",x"c2",x"9c",x"c3"),
  2549 => (x"87",x"c2",x"c1",x"05"),
  2550 => (x"c9",x"49",x"66",x"c4"),
  2551 => (x"c4",x"1e",x"71",x"31"),
  2552 => (x"92",x"d4",x"4a",x"66"),
  2553 => (x"49",x"d9",x"f8",x"c2"),
  2554 => (x"c7",x"fe",x"81",x"72"),
  2555 => (x"49",x"d8",x"87",x"e4"),
  2556 => (x"87",x"dd",x"d5",x"ff"),
  2557 => (x"c2",x"1e",x"c0",x"c8"),
  2558 => (x"fd",x"49",x"f6",x"e6"),
  2559 => (x"ff",x"87",x"df",x"e3"),
  2560 => (x"e0",x"c0",x"48",x"d0"),
  2561 => (x"f6",x"e6",x"c2",x"78"),
  2562 => (x"4a",x"66",x"cc",x"1e"),
  2563 => (x"f8",x"c2",x"92",x"d4"),
  2564 => (x"81",x"72",x"49",x"d9"),
  2565 => (x"87",x"eb",x"c5",x"fe"),
  2566 => (x"ac",x"c1",x"86",x"cc"),
  2567 => (x"87",x"c2",x"c1",x"05"),
  2568 => (x"c9",x"49",x"66",x"c4"),
  2569 => (x"c4",x"1e",x"71",x"31"),
  2570 => (x"92",x"d4",x"4a",x"66"),
  2571 => (x"49",x"d9",x"f8",x"c2"),
  2572 => (x"c6",x"fe",x"81",x"72"),
  2573 => (x"e6",x"c2",x"87",x"dc"),
  2574 => (x"66",x"c8",x"1e",x"f6"),
  2575 => (x"c2",x"92",x"d4",x"4a"),
  2576 => (x"72",x"49",x"d9",x"f8"),
  2577 => (x"eb",x"c3",x"fe",x"81"),
  2578 => (x"ff",x"49",x"d7",x"87"),
  2579 => (x"c8",x"87",x"c2",x"d4"),
  2580 => (x"e6",x"c2",x"1e",x"c0"),
  2581 => (x"e1",x"fd",x"49",x"f6"),
  2582 => (x"86",x"cc",x"87",x"dd"),
  2583 => (x"c0",x"48",x"d0",x"ff"),
  2584 => (x"8e",x"f8",x"78",x"e0"),
  2585 => (x"0e",x"87",x"e7",x"fc"),
  2586 => (x"5d",x"5c",x"5b",x"5e"),
  2587 => (x"4d",x"71",x"1e",x"0e"),
  2588 => (x"d4",x"4c",x"d4",x"ff"),
  2589 => (x"c3",x"48",x"7e",x"66"),
  2590 => (x"c5",x"06",x"a8",x"b7"),
  2591 => (x"c1",x"48",x"c0",x"87"),
  2592 => (x"49",x"75",x"87",x"e2"),
  2593 => (x"87",x"d7",x"d4",x"fe"),
  2594 => (x"66",x"c4",x"1e",x"75"),
  2595 => (x"c2",x"93",x"d4",x"4b"),
  2596 => (x"73",x"83",x"d9",x"f8"),
  2597 => (x"e7",x"fd",x"fd",x"49"),
  2598 => (x"6b",x"83",x"c8",x"87"),
  2599 => (x"48",x"d0",x"ff",x"4b"),
  2600 => (x"dd",x"78",x"e1",x"c8"),
  2601 => (x"c3",x"49",x"73",x"7c"),
  2602 => (x"7c",x"71",x"99",x"ff"),
  2603 => (x"b7",x"c8",x"49",x"73"),
  2604 => (x"99",x"ff",x"c3",x"29"),
  2605 => (x"49",x"73",x"7c",x"71"),
  2606 => (x"c3",x"29",x"b7",x"d0"),
  2607 => (x"7c",x"71",x"99",x"ff"),
  2608 => (x"b7",x"d8",x"49",x"73"),
  2609 => (x"c0",x"7c",x"71",x"29"),
  2610 => (x"7c",x"7c",x"7c",x"7c"),
  2611 => (x"7c",x"7c",x"7c",x"7c"),
  2612 => (x"7c",x"7c",x"7c",x"7c"),
  2613 => (x"c4",x"78",x"e0",x"c0"),
  2614 => (x"49",x"dc",x"1e",x"66"),
  2615 => (x"87",x"d6",x"d2",x"ff"),
  2616 => (x"48",x"73",x"86",x"c8"),
  2617 => (x"87",x"e4",x"fa",x"26"),
  2618 => (x"c4",x"4a",x"71",x"1e"),
  2619 => (x"f7",x"c2",x"49",x"a2"),
  2620 => (x"78",x"6a",x"48",x"f0"),
  2621 => (x"48",x"da",x"db",x"c2"),
  2622 => (x"db",x"c2",x"78",x"69"),
  2623 => (x"e8",x"49",x"bf",x"da"),
  2624 => (x"d3",x"ff",x"87",x"c2"),
  2625 => (x"48",x"c1",x"87",x"ca"),
  2626 => (x"71",x"1e",x"4f",x"26"),
  2627 => (x"49",x"a2",x"c4",x"4a"),
  2628 => (x"bf",x"f0",x"f7",x"c2"),
  2629 => (x"da",x"db",x"c2",x"7a"),
  2630 => (x"4f",x"26",x"79",x"bf"),
  2631 => (x"9a",x"4a",x"71",x"1e"),
  2632 => (x"87",x"ec",x"c0",x"02"),
  2633 => (x"ec",x"f3",x"c2",x"1e"),
  2634 => (x"d3",x"fb",x"fd",x"49"),
  2635 => (x"70",x"86",x"c4",x"87"),
  2636 => (x"87",x"dc",x"02",x"98"),
  2637 => (x"1e",x"f6",x"e6",x"c2"),
  2638 => (x"49",x"ec",x"f3",x"c2"),
  2639 => (x"87",x"f4",x"ff",x"fd"),
  2640 => (x"98",x"70",x"86",x"c4"),
  2641 => (x"c2",x"87",x"c9",x"02"),
  2642 => (x"fe",x"49",x"f6",x"e6"),
  2643 => (x"87",x"c2",x"87",x"da"),
  2644 => (x"4f",x"26",x"48",x"c0"),
  2645 => (x"9a",x"4a",x"71",x"1e"),
  2646 => (x"87",x"ee",x"c0",x"02"),
  2647 => (x"ec",x"f3",x"c2",x"1e"),
  2648 => (x"db",x"fa",x"fd",x"49"),
  2649 => (x"70",x"86",x"c4",x"87"),
  2650 => (x"87",x"de",x"02",x"98"),
  2651 => (x"49",x"f6",x"e6",x"c2"),
  2652 => (x"c2",x"87",x"d7",x"fe"),
  2653 => (x"c2",x"1e",x"f6",x"e6"),
  2654 => (x"fe",x"49",x"ec",x"f3"),
  2655 => (x"c4",x"87",x"c4",x"c0"),
  2656 => (x"02",x"98",x"70",x"86"),
  2657 => (x"48",x"c1",x"87",x"c4"),
  2658 => (x"48",x"c0",x"87",x"c2"),
  2659 => (x"48",x"c0",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

