
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"3e",x"1c",x"00",x"00"),
     1 => (x"00",x"00",x"41",x"63"),
     2 => (x"63",x"41",x"00",x"00"),
     3 => (x"00",x"00",x"1c",x"3e"),
     4 => (x"1c",x"3e",x"2a",x"08"),
     5 => (x"08",x"2a",x"3e",x"1c"),
     6 => (x"3e",x"08",x"08",x"00"),
     7 => (x"00",x"08",x"08",x"3e"),
     8 => (x"e0",x"80",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"60"),
    10 => (x"08",x"08",x"08",x"00"),
    11 => (x"00",x"08",x"08",x"08"),
    12 => (x"60",x"00",x"00",x"00"),
    13 => (x"00",x"00",x"00",x"60"),
    14 => (x"18",x"30",x"60",x"40"),
    15 => (x"01",x"03",x"06",x"0c"),
    16 => (x"59",x"7f",x"3e",x"00"),
    17 => (x"00",x"3e",x"7f",x"4d"),
    18 => (x"7f",x"06",x"04",x"00"),
    19 => (x"00",x"00",x"00",x"7f"),
    20 => (x"71",x"63",x"42",x"00"),
    21 => (x"00",x"46",x"4f",x"59"),
    22 => (x"49",x"63",x"22",x"00"),
    23 => (x"00",x"36",x"7f",x"49"),
    24 => (x"13",x"16",x"1c",x"18"),
    25 => (x"00",x"10",x"7f",x"7f"),
    26 => (x"45",x"67",x"27",x"00"),
    27 => (x"00",x"39",x"7d",x"45"),
    28 => (x"4b",x"7e",x"3c",x"00"),
    29 => (x"00",x"30",x"79",x"49"),
    30 => (x"71",x"01",x"01",x"00"),
    31 => (x"00",x"07",x"0f",x"79"),
    32 => (x"49",x"7f",x"36",x"00"),
    33 => (x"00",x"36",x"7f",x"49"),
    34 => (x"49",x"4f",x"06",x"00"),
    35 => (x"00",x"1e",x"3f",x"69"),
    36 => (x"66",x"00",x"00",x"00"),
    37 => (x"00",x"00",x"00",x"66"),
    38 => (x"e6",x"80",x"00",x"00"),
    39 => (x"00",x"00",x"00",x"66"),
    40 => (x"14",x"08",x"08",x"00"),
    41 => (x"00",x"22",x"22",x"14"),
    42 => (x"14",x"14",x"14",x"00"),
    43 => (x"00",x"14",x"14",x"14"),
    44 => (x"14",x"22",x"22",x"00"),
    45 => (x"00",x"08",x"08",x"14"),
    46 => (x"51",x"03",x"02",x"00"),
    47 => (x"00",x"06",x"0f",x"59"),
    48 => (x"5d",x"41",x"7f",x"3e"),
    49 => (x"00",x"1e",x"1f",x"55"),
    50 => (x"09",x"7f",x"7e",x"00"),
    51 => (x"00",x"7e",x"7f",x"09"),
    52 => (x"49",x"7f",x"7f",x"00"),
    53 => (x"00",x"36",x"7f",x"49"),
    54 => (x"63",x"3e",x"1c",x"00"),
    55 => (x"00",x"41",x"41",x"41"),
    56 => (x"41",x"7f",x"7f",x"00"),
    57 => (x"00",x"1c",x"3e",x"63"),
    58 => (x"49",x"7f",x"7f",x"00"),
    59 => (x"00",x"41",x"41",x"49"),
    60 => (x"09",x"7f",x"7f",x"00"),
    61 => (x"00",x"01",x"01",x"09"),
    62 => (x"41",x"7f",x"3e",x"00"),
    63 => (x"00",x"7a",x"7b",x"49"),
    64 => (x"08",x"7f",x"7f",x"00"),
    65 => (x"00",x"7f",x"7f",x"08"),
    66 => (x"7f",x"41",x"00",x"00"),
    67 => (x"00",x"00",x"41",x"7f"),
    68 => (x"40",x"60",x"20",x"00"),
    69 => (x"00",x"3f",x"7f",x"40"),
    70 => (x"1c",x"08",x"7f",x"7f"),
    71 => (x"00",x"41",x"63",x"36"),
    72 => (x"40",x"7f",x"7f",x"00"),
    73 => (x"00",x"40",x"40",x"40"),
    74 => (x"0c",x"06",x"7f",x"7f"),
    75 => (x"00",x"7f",x"7f",x"06"),
    76 => (x"0c",x"06",x"7f",x"7f"),
    77 => (x"00",x"7f",x"7f",x"18"),
    78 => (x"41",x"7f",x"3e",x"00"),
    79 => (x"00",x"3e",x"7f",x"41"),
    80 => (x"09",x"7f",x"7f",x"00"),
    81 => (x"00",x"06",x"0f",x"09"),
    82 => (x"61",x"41",x"7f",x"3e"),
    83 => (x"00",x"40",x"7e",x"7f"),
    84 => (x"09",x"7f",x"7f",x"00"),
    85 => (x"00",x"66",x"7f",x"19"),
    86 => (x"4d",x"6f",x"26",x"00"),
    87 => (x"00",x"32",x"7b",x"59"),
    88 => (x"7f",x"01",x"01",x"00"),
    89 => (x"00",x"01",x"01",x"7f"),
    90 => (x"40",x"7f",x"3f",x"00"),
    91 => (x"00",x"3f",x"7f",x"40"),
    92 => (x"70",x"3f",x"0f",x"00"),
    93 => (x"00",x"0f",x"3f",x"70"),
    94 => (x"18",x"30",x"7f",x"7f"),
    95 => (x"00",x"7f",x"7f",x"30"),
    96 => (x"1c",x"36",x"63",x"41"),
    97 => (x"41",x"63",x"36",x"1c"),
    98 => (x"7c",x"06",x"03",x"01"),
    99 => (x"01",x"03",x"06",x"7c"),
   100 => (x"4d",x"59",x"71",x"61"),
   101 => (x"00",x"41",x"43",x"47"),
   102 => (x"7f",x"7f",x"00",x"00"),
   103 => (x"00",x"00",x"41",x"41"),
   104 => (x"0c",x"06",x"03",x"01"),
   105 => (x"40",x"60",x"30",x"18"),
   106 => (x"41",x"41",x"00",x"00"),
   107 => (x"00",x"00",x"7f",x"7f"),
   108 => (x"03",x"06",x"0c",x"08"),
   109 => (x"00",x"08",x"0c",x"06"),
   110 => (x"80",x"80",x"80",x"80"),
   111 => (x"00",x"80",x"80",x"80"),
   112 => (x"03",x"00",x"00",x"00"),
   113 => (x"00",x"00",x"04",x"07"),
   114 => (x"54",x"74",x"20",x"00"),
   115 => (x"00",x"78",x"7c",x"54"),
   116 => (x"44",x"7f",x"7f",x"00"),
   117 => (x"00",x"38",x"7c",x"44"),
   118 => (x"44",x"7c",x"38",x"00"),
   119 => (x"00",x"00",x"44",x"44"),
   120 => (x"44",x"7c",x"38",x"00"),
   121 => (x"00",x"7f",x"7f",x"44"),
   122 => (x"54",x"7c",x"38",x"00"),
   123 => (x"00",x"18",x"5c",x"54"),
   124 => (x"7f",x"7e",x"04",x"00"),
   125 => (x"00",x"00",x"05",x"05"),
   126 => (x"a4",x"bc",x"18",x"00"),
   127 => (x"00",x"7c",x"fc",x"a4"),
   128 => (x"04",x"7f",x"7f",x"00"),
   129 => (x"00",x"78",x"7c",x"04"),
   130 => (x"3d",x"00",x"00",x"00"),
   131 => (x"00",x"00",x"40",x"7d"),
   132 => (x"80",x"80",x"80",x"00"),
   133 => (x"00",x"00",x"7d",x"fd"),
   134 => (x"10",x"7f",x"7f",x"00"),
   135 => (x"00",x"44",x"6c",x"38"),
   136 => (x"3f",x"00",x"00",x"00"),
   137 => (x"00",x"00",x"40",x"7f"),
   138 => (x"18",x"0c",x"7c",x"7c"),
   139 => (x"00",x"78",x"7c",x"0c"),
   140 => (x"04",x"7c",x"7c",x"00"),
   141 => (x"00",x"78",x"7c",x"04"),
   142 => (x"44",x"7c",x"38",x"00"),
   143 => (x"00",x"38",x"7c",x"44"),
   144 => (x"24",x"fc",x"fc",x"00"),
   145 => (x"00",x"18",x"3c",x"24"),
   146 => (x"24",x"3c",x"18",x"00"),
   147 => (x"00",x"fc",x"fc",x"24"),
   148 => (x"04",x"7c",x"7c",x"00"),
   149 => (x"00",x"08",x"0c",x"04"),
   150 => (x"54",x"5c",x"48",x"00"),
   151 => (x"00",x"20",x"74",x"54"),
   152 => (x"7f",x"3f",x"04",x"00"),
   153 => (x"00",x"00",x"44",x"44"),
   154 => (x"40",x"7c",x"3c",x"00"),
   155 => (x"00",x"7c",x"7c",x"40"),
   156 => (x"60",x"3c",x"1c",x"00"),
   157 => (x"00",x"1c",x"3c",x"60"),
   158 => (x"30",x"60",x"7c",x"3c"),
   159 => (x"00",x"3c",x"7c",x"60"),
   160 => (x"10",x"38",x"6c",x"44"),
   161 => (x"00",x"44",x"6c",x"38"),
   162 => (x"e0",x"bc",x"1c",x"00"),
   163 => (x"00",x"1c",x"3c",x"60"),
   164 => (x"74",x"64",x"44",x"00"),
   165 => (x"00",x"44",x"4c",x"5c"),
   166 => (x"3e",x"08",x"08",x"00"),
   167 => (x"00",x"41",x"41",x"77"),
   168 => (x"7f",x"00",x"00",x"00"),
   169 => (x"00",x"00",x"00",x"7f"),
   170 => (x"77",x"41",x"41",x"00"),
   171 => (x"00",x"08",x"08",x"3e"),
   172 => (x"03",x"01",x"01",x"02"),
   173 => (x"00",x"01",x"02",x"02"),
   174 => (x"7f",x"7f",x"7f",x"7f"),
   175 => (x"00",x"7f",x"7f",x"7f"),
   176 => (x"1c",x"1c",x"08",x"08"),
   177 => (x"7f",x"7f",x"3e",x"3e"),
   178 => (x"3e",x"3e",x"7f",x"7f"),
   179 => (x"08",x"08",x"1c",x"1c"),
   180 => (x"7c",x"18",x"10",x"00"),
   181 => (x"00",x"10",x"18",x"7c"),
   182 => (x"7c",x"30",x"10",x"00"),
   183 => (x"00",x"10",x"30",x"7c"),
   184 => (x"60",x"60",x"30",x"10"),
   185 => (x"00",x"06",x"1e",x"78"),
   186 => (x"18",x"3c",x"66",x"42"),
   187 => (x"00",x"42",x"66",x"3c"),
   188 => (x"c2",x"6a",x"38",x"78"),
   189 => (x"00",x"38",x"6c",x"c6"),
   190 => (x"60",x"00",x"00",x"60"),
   191 => (x"00",x"60",x"00",x"00"),
   192 => (x"5c",x"5b",x"5e",x"0e"),
   193 => (x"86",x"fc",x"0e",x"5d"),
   194 => (x"f8",x"c2",x"7e",x"71"),
   195 => (x"c0",x"4c",x"bf",x"f8"),
   196 => (x"c4",x"1e",x"c0",x"4b"),
   197 => (x"c4",x"02",x"ab",x"66"),
   198 => (x"c2",x"4d",x"c0",x"87"),
   199 => (x"75",x"4d",x"c1",x"87"),
   200 => (x"ee",x"49",x"73",x"1e"),
   201 => (x"86",x"c8",x"87",x"e3"),
   202 => (x"ef",x"49",x"e0",x"c0"),
   203 => (x"a4",x"c4",x"87",x"ec"),
   204 => (x"f0",x"49",x"6a",x"4a"),
   205 => (x"ca",x"f1",x"87",x"f3"),
   206 => (x"c1",x"84",x"cc",x"87"),
   207 => (x"ab",x"b7",x"c8",x"83"),
   208 => (x"87",x"cd",x"ff",x"04"),
   209 => (x"4d",x"26",x"8e",x"fc"),
   210 => (x"4b",x"26",x"4c",x"26"),
   211 => (x"71",x"1e",x"4f",x"26"),
   212 => (x"fc",x"f8",x"c2",x"4a"),
   213 => (x"fc",x"f8",x"c2",x"5a"),
   214 => (x"49",x"78",x"c7",x"48"),
   215 => (x"26",x"87",x"e1",x"fe"),
   216 => (x"1e",x"73",x"1e",x"4f"),
   217 => (x"b7",x"c0",x"4a",x"71"),
   218 => (x"87",x"d3",x"03",x"aa"),
   219 => (x"bf",x"cc",x"dc",x"c2"),
   220 => (x"c1",x"87",x"c4",x"05"),
   221 => (x"c0",x"87",x"c2",x"4b"),
   222 => (x"d0",x"dc",x"c2",x"4b"),
   223 => (x"c2",x"87",x"c4",x"5b"),
   224 => (x"fc",x"5a",x"d0",x"dc"),
   225 => (x"cc",x"dc",x"c2",x"48"),
   226 => (x"c1",x"4a",x"78",x"bf"),
   227 => (x"a2",x"c0",x"c1",x"9a"),
   228 => (x"87",x"e8",x"ec",x"49"),
   229 => (x"4f",x"26",x"4b",x"26"),
   230 => (x"c4",x"4a",x"71",x"1e"),
   231 => (x"49",x"72",x"1e",x"66"),
   232 => (x"fc",x"87",x"e0",x"eb"),
   233 => (x"1e",x"4f",x"26",x"8e"),
   234 => (x"c3",x"48",x"d4",x"ff"),
   235 => (x"d0",x"ff",x"78",x"ff"),
   236 => (x"78",x"e1",x"c0",x"48"),
   237 => (x"c1",x"48",x"d4",x"ff"),
   238 => (x"c4",x"48",x"71",x"78"),
   239 => (x"08",x"d4",x"ff",x"30"),
   240 => (x"48",x"d0",x"ff",x"78"),
   241 => (x"26",x"78",x"e0",x"c0"),
   242 => (x"5b",x"5e",x"0e",x"4f"),
   243 => (x"f0",x"0e",x"5d",x"5c"),
   244 => (x"c8",x"7e",x"c0",x"86"),
   245 => (x"bf",x"ec",x"48",x"a6"),
   246 => (x"c2",x"80",x"fc",x"78"),
   247 => (x"78",x"bf",x"f8",x"f8"),
   248 => (x"bf",x"c0",x"f9",x"c2"),
   249 => (x"4c",x"bf",x"e8",x"4d"),
   250 => (x"bf",x"cc",x"dc",x"c2"),
   251 => (x"87",x"de",x"e3",x"49"),
   252 => (x"d6",x"e8",x"49",x"c7"),
   253 => (x"c2",x"49",x"70",x"87"),
   254 => (x"87",x"d0",x"05",x"99"),
   255 => (x"bf",x"c4",x"dc",x"c2"),
   256 => (x"c8",x"b9",x"ff",x"49"),
   257 => (x"99",x"c1",x"99",x"66"),
   258 => (x"87",x"c2",x"c2",x"02"),
   259 => (x"cb",x"49",x"e8",x"cf"),
   260 => (x"a6",x"d0",x"87",x"fe"),
   261 => (x"e7",x"49",x"c7",x"58"),
   262 => (x"98",x"70",x"87",x"f1"),
   263 => (x"c8",x"87",x"c9",x"05"),
   264 => (x"99",x"c1",x"49",x"66"),
   265 => (x"87",x"c6",x"c1",x"02"),
   266 => (x"c8",x"4b",x"66",x"cc"),
   267 => (x"bf",x"ec",x"48",x"a6"),
   268 => (x"cc",x"dc",x"c2",x"78"),
   269 => (x"d5",x"e2",x"49",x"bf"),
   270 => (x"cb",x"49",x"73",x"87"),
   271 => (x"98",x"70",x"87",x"de"),
   272 => (x"c2",x"87",x"d7",x"02"),
   273 => (x"49",x"bf",x"c0",x"dc"),
   274 => (x"dc",x"c2",x"b9",x"c1"),
   275 => (x"fd",x"71",x"59",x"c4"),
   276 => (x"e8",x"cf",x"87",x"d5"),
   277 => (x"87",x"f8",x"ca",x"49"),
   278 => (x"49",x"c7",x"4b",x"70"),
   279 => (x"70",x"87",x"ec",x"e6"),
   280 => (x"c6",x"ff",x"05",x"98"),
   281 => (x"49",x"66",x"c8",x"87"),
   282 => (x"fe",x"05",x"99",x"c1"),
   283 => (x"dc",x"c2",x"87",x"fd"),
   284 => (x"c1",x"4a",x"bf",x"cc"),
   285 => (x"d0",x"dc",x"c2",x"ba"),
   286 => (x"7a",x"0a",x"fc",x"5a"),
   287 => (x"c1",x"9a",x"c1",x"0a"),
   288 => (x"e8",x"49",x"a2",x"c0"),
   289 => (x"da",x"c1",x"87",x"f6"),
   290 => (x"87",x"ff",x"e5",x"49"),
   291 => (x"dc",x"c2",x"7e",x"c1"),
   292 => (x"66",x"c8",x"48",x"c4"),
   293 => (x"cc",x"dc",x"c2",x"78"),
   294 => (x"c7",x"c1",x"05",x"bf"),
   295 => (x"c0",x"c0",x"c8",x"87"),
   296 => (x"f0",x"db",x"c2",x"4b"),
   297 => (x"49",x"15",x"4d",x"7e"),
   298 => (x"87",x"df",x"e5",x"49"),
   299 => (x"c0",x"02",x"98",x"70"),
   300 => (x"b4",x"73",x"87",x"c2"),
   301 => (x"05",x"2b",x"b7",x"c1"),
   302 => (x"74",x"87",x"eb",x"ff"),
   303 => (x"99",x"ff",x"c3",x"49"),
   304 => (x"49",x"c0",x"1e",x"71"),
   305 => (x"74",x"87",x"d1",x"fb"),
   306 => (x"29",x"b7",x"c8",x"49"),
   307 => (x"49",x"c1",x"1e",x"71"),
   308 => (x"c8",x"87",x"c5",x"fb"),
   309 => (x"49",x"fd",x"c3",x"86"),
   310 => (x"c3",x"87",x"f0",x"e4"),
   311 => (x"ea",x"e4",x"49",x"fa"),
   312 => (x"87",x"fe",x"c7",x"87"),
   313 => (x"ff",x"c3",x"49",x"74"),
   314 => (x"2c",x"b7",x"c8",x"99"),
   315 => (x"9c",x"74",x"b4",x"71"),
   316 => (x"87",x"e5",x"c0",x"02"),
   317 => (x"ff",x"48",x"a6",x"c8"),
   318 => (x"c8",x"78",x"bf",x"c8"),
   319 => (x"dc",x"c2",x"49",x"66"),
   320 => (x"c2",x"89",x"bf",x"c8"),
   321 => (x"c0",x"03",x"a9",x"e0"),
   322 => (x"4c",x"c0",x"87",x"c5"),
   323 => (x"c2",x"87",x"d0",x"c0"),
   324 => (x"c8",x"48",x"c8",x"dc"),
   325 => (x"c6",x"c0",x"78",x"66"),
   326 => (x"c8",x"dc",x"c2",x"87"),
   327 => (x"74",x"78",x"c0",x"48"),
   328 => (x"05",x"99",x"c8",x"49"),
   329 => (x"c3",x"87",x"ce",x"c0"),
   330 => (x"de",x"e3",x"49",x"f5"),
   331 => (x"c2",x"49",x"70",x"87"),
   332 => (x"e7",x"c0",x"02",x"99"),
   333 => (x"fc",x"f8",x"c2",x"87"),
   334 => (x"ca",x"c0",x"02",x"bf"),
   335 => (x"88",x"c1",x"48",x"87"),
   336 => (x"58",x"c0",x"f9",x"c2"),
   337 => (x"c4",x"87",x"d3",x"c0"),
   338 => (x"e0",x"c1",x"48",x"66"),
   339 => (x"6e",x"7e",x"70",x"80"),
   340 => (x"c5",x"c0",x"02",x"bf"),
   341 => (x"49",x"ff",x"4b",x"87"),
   342 => (x"7e",x"c1",x"0f",x"73"),
   343 => (x"99",x"c4",x"49",x"74"),
   344 => (x"87",x"ce",x"c0",x"05"),
   345 => (x"e2",x"49",x"f2",x"c3"),
   346 => (x"49",x"70",x"87",x"e1"),
   347 => (x"c0",x"02",x"99",x"c2"),
   348 => (x"f8",x"c2",x"87",x"ed"),
   349 => (x"48",x"7e",x"bf",x"fc"),
   350 => (x"03",x"a8",x"b7",x"c7"),
   351 => (x"6e",x"87",x"cb",x"c0"),
   352 => (x"c2",x"80",x"c1",x"48"),
   353 => (x"c0",x"58",x"c0",x"f9"),
   354 => (x"66",x"c4",x"87",x"d3"),
   355 => (x"80",x"e0",x"c1",x"48"),
   356 => (x"bf",x"6e",x"7e",x"70"),
   357 => (x"87",x"c5",x"c0",x"02"),
   358 => (x"73",x"49",x"fe",x"4b"),
   359 => (x"c3",x"7e",x"c1",x"0f"),
   360 => (x"e6",x"e1",x"49",x"fd"),
   361 => (x"c2",x"49",x"70",x"87"),
   362 => (x"e3",x"c0",x"02",x"99"),
   363 => (x"fc",x"f8",x"c2",x"87"),
   364 => (x"c9",x"c0",x"02",x"bf"),
   365 => (x"fc",x"f8",x"c2",x"87"),
   366 => (x"c0",x"78",x"c0",x"48"),
   367 => (x"66",x"c4",x"87",x"d0"),
   368 => (x"82",x"e0",x"c1",x"4a"),
   369 => (x"c5",x"c0",x"02",x"6a"),
   370 => (x"49",x"fd",x"4b",x"87"),
   371 => (x"7e",x"c1",x"0f",x"73"),
   372 => (x"e0",x"49",x"fa",x"c3"),
   373 => (x"49",x"70",x"87",x"f5"),
   374 => (x"c0",x"02",x"99",x"c2"),
   375 => (x"f8",x"c2",x"87",x"ea"),
   376 => (x"c7",x"48",x"bf",x"fc"),
   377 => (x"c0",x"03",x"a8",x"b7"),
   378 => (x"f8",x"c2",x"87",x"c9"),
   379 => (x"78",x"c7",x"48",x"fc"),
   380 => (x"c4",x"87",x"d3",x"c0"),
   381 => (x"e0",x"c1",x"48",x"66"),
   382 => (x"6e",x"7e",x"70",x"80"),
   383 => (x"c5",x"c0",x"02",x"bf"),
   384 => (x"49",x"fc",x"4b",x"87"),
   385 => (x"7e",x"c1",x"0f",x"73"),
   386 => (x"f0",x"c3",x"48",x"74"),
   387 => (x"58",x"a6",x"cc",x"98"),
   388 => (x"c0",x"05",x"98",x"70"),
   389 => (x"da",x"c1",x"87",x"cf"),
   390 => (x"ee",x"df",x"ff",x"49"),
   391 => (x"c2",x"49",x"70",x"87"),
   392 => (x"c1",x"c2",x"02",x"99"),
   393 => (x"49",x"e8",x"cf",x"87"),
   394 => (x"d0",x"87",x"e5",x"c3"),
   395 => (x"f8",x"c2",x"58",x"a6"),
   396 => (x"50",x"c0",x"48",x"f4"),
   397 => (x"97",x"f4",x"f8",x"c2"),
   398 => (x"d9",x"c1",x"05",x"bf"),
   399 => (x"05",x"66",x"c8",x"87"),
   400 => (x"c1",x"87",x"cd",x"c0"),
   401 => (x"df",x"ff",x"49",x"da"),
   402 => (x"98",x"70",x"87",x"c1"),
   403 => (x"87",x"c6",x"c1",x"02"),
   404 => (x"49",x"4b",x"bf",x"e8"),
   405 => (x"c8",x"99",x"ff",x"c3"),
   406 => (x"b3",x"71",x"2b",x"b7"),
   407 => (x"bf",x"cc",x"dc",x"c2"),
   408 => (x"e9",x"d9",x"ff",x"49"),
   409 => (x"49",x"66",x"cc",x"87"),
   410 => (x"70",x"87",x"f1",x"c2"),
   411 => (x"c6",x"c0",x"02",x"98"),
   412 => (x"f4",x"f8",x"c2",x"87"),
   413 => (x"c2",x"50",x"c1",x"48"),
   414 => (x"bf",x"97",x"f4",x"f8"),
   415 => (x"87",x"d6",x"c0",x"05"),
   416 => (x"f0",x"c3",x"49",x"73"),
   417 => (x"c7",x"ff",x"05",x"99"),
   418 => (x"49",x"da",x"c1",x"87"),
   419 => (x"87",x"fb",x"dd",x"ff"),
   420 => (x"fe",x"05",x"98",x"70"),
   421 => (x"f8",x"c2",x"87",x"fa"),
   422 => (x"4b",x"49",x"bf",x"fc"),
   423 => (x"66",x"c4",x"93",x"cc"),
   424 => (x"71",x"4b",x"6b",x"83"),
   425 => (x"9d",x"75",x"0f",x"73"),
   426 => (x"87",x"e9",x"c0",x"02"),
   427 => (x"e4",x"c0",x"02",x"6d"),
   428 => (x"ff",x"49",x"6d",x"87"),
   429 => (x"70",x"87",x"d4",x"dd"),
   430 => (x"02",x"99",x"c1",x"49"),
   431 => (x"c4",x"87",x"cb",x"c0"),
   432 => (x"f8",x"c2",x"4b",x"a5"),
   433 => (x"6b",x"49",x"bf",x"fc"),
   434 => (x"85",x"c8",x"0f",x"4b"),
   435 => (x"87",x"c5",x"c0",x"02"),
   436 => (x"dc",x"ff",x"05",x"6d"),
   437 => (x"c0",x"02",x"6e",x"87"),
   438 => (x"f8",x"c2",x"87",x"c8"),
   439 => (x"f0",x"49",x"bf",x"fc"),
   440 => (x"8e",x"f0",x"87",x"de"),
   441 => (x"4c",x"26",x"4d",x"26"),
   442 => (x"4f",x"26",x"4b",x"26"),
   443 => (x"00",x"00",x"00",x"10"),
   444 => (x"14",x"11",x"12",x"58"),
   445 => (x"23",x"1c",x"1b",x"1d"),
   446 => (x"94",x"91",x"59",x"5a"),
   447 => (x"f4",x"eb",x"f2",x"f5"),
   448 => (x"00",x"00",x"00",x"00"),
   449 => (x"00",x"00",x"00",x"00"),
   450 => (x"00",x"00",x"00",x"00"),
   451 => (x"00",x"00",x"00",x"00"),
   452 => (x"ff",x"4a",x"71",x"1e"),
   453 => (x"72",x"49",x"bf",x"c8"),
   454 => (x"4f",x"26",x"48",x"a1"),
   455 => (x"bf",x"c8",x"ff",x"1e"),
   456 => (x"c0",x"c0",x"fe",x"89"),
   457 => (x"a9",x"c0",x"c0",x"c0"),
   458 => (x"c0",x"87",x"c4",x"01"),
   459 => (x"c1",x"87",x"c2",x"4a"),
   460 => (x"26",x"48",x"72",x"4a"),
   461 => (x"5b",x"5e",x"0e",x"4f"),
   462 => (x"71",x"0e",x"5d",x"5c"),
   463 => (x"4c",x"d4",x"ff",x"4b"),
   464 => (x"c0",x"48",x"66",x"d0"),
   465 => (x"ff",x"49",x"d6",x"78"),
   466 => (x"c3",x"87",x"fd",x"db"),
   467 => (x"49",x"6c",x"7c",x"ff"),
   468 => (x"71",x"99",x"ff",x"c3"),
   469 => (x"f0",x"c3",x"49",x"4d"),
   470 => (x"a9",x"e0",x"c1",x"99"),
   471 => (x"c3",x"87",x"cb",x"05"),
   472 => (x"48",x"6c",x"7c",x"ff"),
   473 => (x"66",x"d0",x"98",x"c3"),
   474 => (x"ff",x"c3",x"78",x"08"),
   475 => (x"49",x"4a",x"6c",x"7c"),
   476 => (x"ff",x"c3",x"31",x"c8"),
   477 => (x"71",x"4a",x"6c",x"7c"),
   478 => (x"c8",x"49",x"72",x"b2"),
   479 => (x"7c",x"ff",x"c3",x"31"),
   480 => (x"b2",x"71",x"4a",x"6c"),
   481 => (x"31",x"c8",x"49",x"72"),
   482 => (x"6c",x"7c",x"ff",x"c3"),
   483 => (x"ff",x"b2",x"71",x"4a"),
   484 => (x"e0",x"c0",x"48",x"d0"),
   485 => (x"02",x"9b",x"73",x"78"),
   486 => (x"7b",x"72",x"87",x"c2"),
   487 => (x"4d",x"26",x"48",x"75"),
   488 => (x"4b",x"26",x"4c",x"26"),
   489 => (x"26",x"1e",x"4f",x"26"),
   490 => (x"5b",x"5e",x"0e",x"4f"),
   491 => (x"86",x"f8",x"0e",x"5c"),
   492 => (x"a6",x"c8",x"1e",x"76"),
   493 => (x"87",x"fd",x"fd",x"49"),
   494 => (x"4b",x"70",x"86",x"c4"),
   495 => (x"a8",x"c4",x"48",x"6e"),
   496 => (x"87",x"fb",x"c2",x"03"),
   497 => (x"f0",x"c3",x"4a",x"73"),
   498 => (x"aa",x"d0",x"c1",x"9a"),
   499 => (x"c1",x"87",x"c7",x"02"),
   500 => (x"c2",x"05",x"aa",x"e0"),
   501 => (x"49",x"73",x"87",x"e9"),
   502 => (x"c3",x"02",x"99",x"c8"),
   503 => (x"87",x"c6",x"ff",x"87"),
   504 => (x"9c",x"c3",x"4c",x"73"),
   505 => (x"c1",x"05",x"ac",x"c2"),
   506 => (x"66",x"c4",x"87",x"c4"),
   507 => (x"71",x"31",x"c9",x"49"),
   508 => (x"4a",x"66",x"c4",x"1e"),
   509 => (x"c2",x"92",x"cc",x"c1"),
   510 => (x"72",x"49",x"c4",x"f9"),
   511 => (x"e9",x"cb",x"fe",x"81"),
   512 => (x"ff",x"49",x"d8",x"87"),
   513 => (x"c8",x"87",x"c1",x"d9"),
   514 => (x"e5",x"c2",x"1e",x"c0"),
   515 => (x"e5",x"fd",x"49",x"fc"),
   516 => (x"d0",x"ff",x"87",x"c4"),
   517 => (x"78",x"e0",x"c0",x"48"),
   518 => (x"1e",x"fc",x"e5",x"c2"),
   519 => (x"c1",x"4a",x"66",x"cc"),
   520 => (x"f9",x"c2",x"92",x"cc"),
   521 => (x"81",x"72",x"49",x"c4"),
   522 => (x"87",x"ff",x"c9",x"fe"),
   523 => (x"ac",x"c1",x"86",x"cc"),
   524 => (x"87",x"cb",x"c1",x"05"),
   525 => (x"fd",x"49",x"ee",x"c0"),
   526 => (x"c4",x"87",x"d1",x"e1"),
   527 => (x"31",x"c9",x"49",x"66"),
   528 => (x"66",x"c4",x"1e",x"71"),
   529 => (x"92",x"cc",x"c1",x"4a"),
   530 => (x"49",x"c4",x"f9",x"c2"),
   531 => (x"ca",x"fe",x"81",x"72"),
   532 => (x"e5",x"c2",x"87",x"d8"),
   533 => (x"66",x"c8",x"1e",x"fc"),
   534 => (x"92",x"cc",x"c1",x"4a"),
   535 => (x"49",x"c4",x"f9",x"c2"),
   536 => (x"c8",x"fe",x"81",x"72"),
   537 => (x"49",x"d7",x"87",x"c6"),
   538 => (x"87",x"dc",x"d7",x"ff"),
   539 => (x"c2",x"1e",x"c0",x"c8"),
   540 => (x"fd",x"49",x"fc",x"e5"),
   541 => (x"cc",x"87",x"fc",x"e2"),
   542 => (x"48",x"d0",x"ff",x"86"),
   543 => (x"f8",x"78",x"e0",x"c0"),
   544 => (x"26",x"4c",x"26",x"8e"),
   545 => (x"1e",x"4f",x"26",x"4b"),
   546 => (x"b7",x"c4",x"4a",x"71"),
   547 => (x"87",x"ce",x"03",x"aa"),
   548 => (x"cc",x"c1",x"49",x"72"),
   549 => (x"c4",x"f9",x"c2",x"91"),
   550 => (x"81",x"c8",x"c1",x"81"),
   551 => (x"4f",x"26",x"79",x"c0"),
   552 => (x"5c",x"5b",x"5e",x"0e"),
   553 => (x"86",x"fc",x"0e",x"5d"),
   554 => (x"d4",x"ff",x"4a",x"71"),
   555 => (x"d4",x"4c",x"c0",x"4b"),
   556 => (x"b7",x"c3",x"4d",x"66"),
   557 => (x"c2",x"c2",x"01",x"ad"),
   558 => (x"02",x"9a",x"72",x"87"),
   559 => (x"1e",x"87",x"ec",x"c0"),
   560 => (x"cc",x"c1",x"49",x"75"),
   561 => (x"c4",x"f9",x"c2",x"91"),
   562 => (x"c8",x"80",x"71",x"48"),
   563 => (x"66",x"c4",x"58",x"a6"),
   564 => (x"e3",x"c1",x"fe",x"49"),
   565 => (x"70",x"86",x"c4",x"87"),
   566 => (x"87",x"d4",x"02",x"98"),
   567 => (x"c8",x"c1",x"49",x"6e"),
   568 => (x"6e",x"79",x"c1",x"81"),
   569 => (x"69",x"81",x"c8",x"49"),
   570 => (x"75",x"87",x"c5",x"4c"),
   571 => (x"87",x"d7",x"fe",x"49"),
   572 => (x"c8",x"48",x"d0",x"ff"),
   573 => (x"7b",x"dd",x"78",x"e1"),
   574 => (x"ff",x"c3",x"48",x"74"),
   575 => (x"74",x"7b",x"70",x"98"),
   576 => (x"29",x"b7",x"c8",x"49"),
   577 => (x"ff",x"c3",x"48",x"71"),
   578 => (x"74",x"7b",x"70",x"98"),
   579 => (x"29",x"b7",x"d0",x"49"),
   580 => (x"ff",x"c3",x"48",x"71"),
   581 => (x"74",x"7b",x"70",x"98"),
   582 => (x"28",x"b7",x"d8",x"48"),
   583 => (x"7b",x"c0",x"7b",x"70"),
   584 => (x"7b",x"7b",x"7b",x"7b"),
   585 => (x"7b",x"7b",x"7b",x"7b"),
   586 => (x"ff",x"7b",x"7b",x"7b"),
   587 => (x"e0",x"c0",x"48",x"d0"),
   588 => (x"dc",x"1e",x"75",x"78"),
   589 => (x"f4",x"d4",x"ff",x"49"),
   590 => (x"fc",x"86",x"c4",x"87"),
   591 => (x"26",x"4d",x"26",x"8e"),
   592 => (x"26",x"4b",x"26",x"4c"),
   593 => (x"00",x"1b",x"f3",x"4f"),
   594 => (x"00",x"1b",x"f3",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

