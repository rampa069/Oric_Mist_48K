
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"14",x"22",x"22",x"00"),
     1 => (x"00",x"08",x"08",x"14"),
     2 => (x"51",x"03",x"02",x"00"),
     3 => (x"00",x"06",x"0f",x"59"),
     4 => (x"5d",x"41",x"7f",x"3e"),
     5 => (x"00",x"1e",x"1f",x"55"),
     6 => (x"09",x"7f",x"7e",x"00"),
     7 => (x"00",x"7e",x"7f",x"09"),
     8 => (x"49",x"7f",x"7f",x"00"),
     9 => (x"00",x"36",x"7f",x"49"),
    10 => (x"63",x"3e",x"1c",x"00"),
    11 => (x"00",x"41",x"41",x"41"),
    12 => (x"41",x"7f",x"7f",x"00"),
    13 => (x"00",x"1c",x"3e",x"63"),
    14 => (x"49",x"7f",x"7f",x"00"),
    15 => (x"00",x"41",x"41",x"49"),
    16 => (x"09",x"7f",x"7f",x"00"),
    17 => (x"00",x"01",x"01",x"09"),
    18 => (x"41",x"7f",x"3e",x"00"),
    19 => (x"00",x"7a",x"7b",x"49"),
    20 => (x"08",x"7f",x"7f",x"00"),
    21 => (x"00",x"7f",x"7f",x"08"),
    22 => (x"7f",x"41",x"00",x"00"),
    23 => (x"00",x"00",x"41",x"7f"),
    24 => (x"40",x"60",x"20",x"00"),
    25 => (x"00",x"3f",x"7f",x"40"),
    26 => (x"1c",x"08",x"7f",x"7f"),
    27 => (x"00",x"41",x"63",x"36"),
    28 => (x"40",x"7f",x"7f",x"00"),
    29 => (x"00",x"40",x"40",x"40"),
    30 => (x"0c",x"06",x"7f",x"7f"),
    31 => (x"00",x"7f",x"7f",x"06"),
    32 => (x"0c",x"06",x"7f",x"7f"),
    33 => (x"00",x"7f",x"7f",x"18"),
    34 => (x"41",x"7f",x"3e",x"00"),
    35 => (x"00",x"3e",x"7f",x"41"),
    36 => (x"09",x"7f",x"7f",x"00"),
    37 => (x"00",x"06",x"0f",x"09"),
    38 => (x"61",x"41",x"7f",x"3e"),
    39 => (x"00",x"40",x"7e",x"7f"),
    40 => (x"09",x"7f",x"7f",x"00"),
    41 => (x"00",x"66",x"7f",x"19"),
    42 => (x"4d",x"6f",x"26",x"00"),
    43 => (x"00",x"32",x"7b",x"59"),
    44 => (x"7f",x"01",x"01",x"00"),
    45 => (x"00",x"01",x"01",x"7f"),
    46 => (x"40",x"7f",x"3f",x"00"),
    47 => (x"00",x"3f",x"7f",x"40"),
    48 => (x"70",x"3f",x"0f",x"00"),
    49 => (x"00",x"0f",x"3f",x"70"),
    50 => (x"18",x"30",x"7f",x"7f"),
    51 => (x"00",x"7f",x"7f",x"30"),
    52 => (x"1c",x"36",x"63",x"41"),
    53 => (x"41",x"63",x"36",x"1c"),
    54 => (x"7c",x"06",x"03",x"01"),
    55 => (x"01",x"03",x"06",x"7c"),
    56 => (x"4d",x"59",x"71",x"61"),
    57 => (x"00",x"41",x"43",x"47"),
    58 => (x"7f",x"7f",x"00",x"00"),
    59 => (x"00",x"00",x"41",x"41"),
    60 => (x"0c",x"06",x"03",x"01"),
    61 => (x"40",x"60",x"30",x"18"),
    62 => (x"41",x"41",x"00",x"00"),
    63 => (x"00",x"00",x"7f",x"7f"),
    64 => (x"03",x"06",x"0c",x"08"),
    65 => (x"00",x"08",x"0c",x"06"),
    66 => (x"80",x"80",x"80",x"80"),
    67 => (x"00",x"80",x"80",x"80"),
    68 => (x"03",x"00",x"00",x"00"),
    69 => (x"00",x"00",x"04",x"07"),
    70 => (x"54",x"74",x"20",x"00"),
    71 => (x"00",x"78",x"7c",x"54"),
    72 => (x"44",x"7f",x"7f",x"00"),
    73 => (x"00",x"38",x"7c",x"44"),
    74 => (x"44",x"7c",x"38",x"00"),
    75 => (x"00",x"00",x"44",x"44"),
    76 => (x"44",x"7c",x"38",x"00"),
    77 => (x"00",x"7f",x"7f",x"44"),
    78 => (x"54",x"7c",x"38",x"00"),
    79 => (x"00",x"18",x"5c",x"54"),
    80 => (x"7f",x"7e",x"04",x"00"),
    81 => (x"00",x"00",x"05",x"05"),
    82 => (x"a4",x"bc",x"18",x"00"),
    83 => (x"00",x"7c",x"fc",x"a4"),
    84 => (x"04",x"7f",x"7f",x"00"),
    85 => (x"00",x"78",x"7c",x"04"),
    86 => (x"3d",x"00",x"00",x"00"),
    87 => (x"00",x"00",x"40",x"7d"),
    88 => (x"80",x"80",x"80",x"00"),
    89 => (x"00",x"00",x"7d",x"fd"),
    90 => (x"10",x"7f",x"7f",x"00"),
    91 => (x"00",x"44",x"6c",x"38"),
    92 => (x"3f",x"00",x"00",x"00"),
    93 => (x"00",x"00",x"40",x"7f"),
    94 => (x"18",x"0c",x"7c",x"7c"),
    95 => (x"00",x"78",x"7c",x"0c"),
    96 => (x"04",x"7c",x"7c",x"00"),
    97 => (x"00",x"78",x"7c",x"04"),
    98 => (x"44",x"7c",x"38",x"00"),
    99 => (x"00",x"38",x"7c",x"44"),
   100 => (x"24",x"fc",x"fc",x"00"),
   101 => (x"00",x"18",x"3c",x"24"),
   102 => (x"24",x"3c",x"18",x"00"),
   103 => (x"00",x"fc",x"fc",x"24"),
   104 => (x"04",x"7c",x"7c",x"00"),
   105 => (x"00",x"08",x"0c",x"04"),
   106 => (x"54",x"5c",x"48",x"00"),
   107 => (x"00",x"20",x"74",x"54"),
   108 => (x"7f",x"3f",x"04",x"00"),
   109 => (x"00",x"00",x"44",x"44"),
   110 => (x"40",x"7c",x"3c",x"00"),
   111 => (x"00",x"7c",x"7c",x"40"),
   112 => (x"60",x"3c",x"1c",x"00"),
   113 => (x"00",x"1c",x"3c",x"60"),
   114 => (x"30",x"60",x"7c",x"3c"),
   115 => (x"00",x"3c",x"7c",x"60"),
   116 => (x"10",x"38",x"6c",x"44"),
   117 => (x"00",x"44",x"6c",x"38"),
   118 => (x"e0",x"bc",x"1c",x"00"),
   119 => (x"00",x"1c",x"3c",x"60"),
   120 => (x"74",x"64",x"44",x"00"),
   121 => (x"00",x"44",x"4c",x"5c"),
   122 => (x"3e",x"08",x"08",x"00"),
   123 => (x"00",x"41",x"41",x"77"),
   124 => (x"7f",x"00",x"00",x"00"),
   125 => (x"00",x"00",x"00",x"7f"),
   126 => (x"77",x"41",x"41",x"00"),
   127 => (x"00",x"08",x"08",x"3e"),
   128 => (x"03",x"01",x"01",x"02"),
   129 => (x"00",x"01",x"02",x"02"),
   130 => (x"7f",x"7f",x"7f",x"7f"),
   131 => (x"00",x"7f",x"7f",x"7f"),
   132 => (x"1c",x"1c",x"08",x"08"),
   133 => (x"7f",x"7f",x"3e",x"3e"),
   134 => (x"3e",x"3e",x"7f",x"7f"),
   135 => (x"08",x"08",x"1c",x"1c"),
   136 => (x"7c",x"18",x"10",x"00"),
   137 => (x"00",x"10",x"18",x"7c"),
   138 => (x"7c",x"30",x"10",x"00"),
   139 => (x"00",x"10",x"30",x"7c"),
   140 => (x"60",x"60",x"30",x"10"),
   141 => (x"00",x"06",x"1e",x"78"),
   142 => (x"18",x"3c",x"66",x"42"),
   143 => (x"00",x"42",x"66",x"3c"),
   144 => (x"c2",x"6a",x"38",x"78"),
   145 => (x"00",x"38",x"6c",x"c6"),
   146 => (x"60",x"00",x"00",x"60"),
   147 => (x"00",x"60",x"00",x"00"),
   148 => (x"5c",x"5b",x"5e",x"0e"),
   149 => (x"71",x"1e",x"0e",x"5d"),
   150 => (x"d1",x"f8",x"c2",x"4c"),
   151 => (x"4b",x"c0",x"4d",x"bf"),
   152 => (x"ab",x"74",x"1e",x"c0"),
   153 => (x"c4",x"87",x"c7",x"02"),
   154 => (x"78",x"c0",x"48",x"a6"),
   155 => (x"a6",x"c4",x"87",x"c5"),
   156 => (x"c4",x"78",x"c1",x"48"),
   157 => (x"49",x"73",x"1e",x"66"),
   158 => (x"c8",x"87",x"df",x"ee"),
   159 => (x"49",x"e0",x"c0",x"86"),
   160 => (x"c4",x"87",x"ef",x"ef"),
   161 => (x"49",x"6a",x"4a",x"a5"),
   162 => (x"f1",x"87",x"f0",x"f0"),
   163 => (x"85",x"cb",x"87",x"c6"),
   164 => (x"b7",x"c8",x"83",x"c1"),
   165 => (x"c7",x"ff",x"04",x"ab"),
   166 => (x"4d",x"26",x"26",x"87"),
   167 => (x"4b",x"26",x"4c",x"26"),
   168 => (x"71",x"1e",x"4f",x"26"),
   169 => (x"d5",x"f8",x"c2",x"4a"),
   170 => (x"d5",x"f8",x"c2",x"5a"),
   171 => (x"49",x"78",x"c7",x"48"),
   172 => (x"26",x"87",x"dd",x"fe"),
   173 => (x"1e",x"73",x"1e",x"4f"),
   174 => (x"b7",x"c0",x"4a",x"71"),
   175 => (x"87",x"d3",x"03",x"aa"),
   176 => (x"bf",x"f6",x"db",x"c2"),
   177 => (x"c1",x"87",x"c4",x"05"),
   178 => (x"c0",x"87",x"c2",x"4b"),
   179 => (x"fa",x"db",x"c2",x"4b"),
   180 => (x"c2",x"87",x"c4",x"5b"),
   181 => (x"c2",x"5a",x"fa",x"db"),
   182 => (x"4a",x"bf",x"f6",x"db"),
   183 => (x"c0",x"c1",x"9a",x"c1"),
   184 => (x"e8",x"ec",x"49",x"a2"),
   185 => (x"de",x"db",x"c2",x"87"),
   186 => (x"db",x"c2",x"49",x"bf"),
   187 => (x"fc",x"b1",x"bf",x"f6"),
   188 => (x"fe",x"78",x"71",x"48"),
   189 => (x"71",x"1e",x"87",x"e8"),
   190 => (x"1e",x"66",x"c4",x"4a"),
   191 => (x"e7",x"ea",x"49",x"72"),
   192 => (x"4f",x"26",x"26",x"87"),
   193 => (x"ff",x"4a",x"71",x"1e"),
   194 => (x"ff",x"c3",x"48",x"d4"),
   195 => (x"48",x"d0",x"ff",x"78"),
   196 => (x"ff",x"78",x"e1",x"c0"),
   197 => (x"78",x"c1",x"48",x"d4"),
   198 => (x"31",x"c4",x"49",x"72"),
   199 => (x"d0",x"ff",x"78",x"71"),
   200 => (x"78",x"e0",x"c0",x"48"),
   201 => (x"c2",x"1e",x"4f",x"26"),
   202 => (x"49",x"bf",x"f6",x"db"),
   203 => (x"c2",x"87",x"ca",x"e6"),
   204 => (x"e8",x"48",x"c9",x"f8"),
   205 => (x"f8",x"c2",x"78",x"bf"),
   206 => (x"bf",x"ec",x"48",x"c5"),
   207 => (x"c9",x"f8",x"c2",x"78"),
   208 => (x"c3",x"49",x"4a",x"bf"),
   209 => (x"b7",x"c8",x"99",x"ff"),
   210 => (x"71",x"48",x"72",x"2a"),
   211 => (x"d1",x"f8",x"c2",x"b0"),
   212 => (x"0e",x"4f",x"26",x"58"),
   213 => (x"5d",x"5c",x"5b",x"5e"),
   214 => (x"ff",x"4b",x"71",x"0e"),
   215 => (x"f8",x"c2",x"87",x"c8"),
   216 => (x"50",x"c0",x"48",x"c4"),
   217 => (x"f0",x"e5",x"49",x"73"),
   218 => (x"4c",x"49",x"70",x"87"),
   219 => (x"ee",x"cb",x"9c",x"c2"),
   220 => (x"87",x"ca",x"ce",x"49"),
   221 => (x"c2",x"4d",x"49",x"70"),
   222 => (x"bf",x"97",x"c4",x"f8"),
   223 => (x"87",x"e2",x"c1",x"05"),
   224 => (x"c2",x"49",x"66",x"d0"),
   225 => (x"99",x"bf",x"cd",x"f8"),
   226 => (x"d4",x"87",x"d6",x"05"),
   227 => (x"f8",x"c2",x"49",x"66"),
   228 => (x"05",x"99",x"bf",x"c5"),
   229 => (x"49",x"73",x"87",x"cb"),
   230 => (x"70",x"87",x"fe",x"e4"),
   231 => (x"c1",x"c1",x"02",x"98"),
   232 => (x"fe",x"4c",x"c1",x"87"),
   233 => (x"49",x"75",x"87",x"c0"),
   234 => (x"70",x"87",x"df",x"cd"),
   235 => (x"87",x"c6",x"02",x"98"),
   236 => (x"48",x"c4",x"f8",x"c2"),
   237 => (x"f8",x"c2",x"50",x"c1"),
   238 => (x"05",x"bf",x"97",x"c4"),
   239 => (x"c2",x"87",x"e3",x"c0"),
   240 => (x"49",x"bf",x"cd",x"f8"),
   241 => (x"05",x"99",x"66",x"d0"),
   242 => (x"c2",x"87",x"d6",x"ff"),
   243 => (x"49",x"bf",x"c5",x"f8"),
   244 => (x"05",x"99",x"66",x"d4"),
   245 => (x"73",x"87",x"ca",x"ff"),
   246 => (x"87",x"fd",x"e3",x"49"),
   247 => (x"fe",x"05",x"98",x"70"),
   248 => (x"48",x"74",x"87",x"ff"),
   249 => (x"0e",x"87",x"f3",x"fa"),
   250 => (x"5d",x"5c",x"5b",x"5e"),
   251 => (x"c0",x"86",x"f4",x"0e"),
   252 => (x"bf",x"ec",x"4c",x"4d"),
   253 => (x"48",x"a6",x"c4",x"7e"),
   254 => (x"bf",x"d1",x"f8",x"c2"),
   255 => (x"1e",x"1e",x"c0",x"78"),
   256 => (x"fd",x"49",x"f7",x"c1"),
   257 => (x"86",x"c8",x"87",x"cd"),
   258 => (x"c0",x"02",x"98",x"70"),
   259 => (x"db",x"c2",x"87",x"f3"),
   260 => (x"c4",x"05",x"bf",x"de"),
   261 => (x"c2",x"7e",x"c1",x"87"),
   262 => (x"c2",x"7e",x"c0",x"87"),
   263 => (x"6e",x"48",x"de",x"db"),
   264 => (x"1e",x"fc",x"ca",x"78"),
   265 => (x"c9",x"02",x"66",x"c4"),
   266 => (x"48",x"a6",x"c4",x"87"),
   267 => (x"78",x"f1",x"d9",x"c2"),
   268 => (x"a6",x"c4",x"87",x"c7"),
   269 => (x"fc",x"d9",x"c2",x"48"),
   270 => (x"49",x"66",x"c4",x"78"),
   271 => (x"c4",x"87",x"c9",x"c9"),
   272 => (x"c0",x"1e",x"c1",x"86"),
   273 => (x"fc",x"49",x"c7",x"1e"),
   274 => (x"86",x"c8",x"87",x"c9"),
   275 => (x"cd",x"02",x"98",x"70"),
   276 => (x"f9",x"49",x"ff",x"87"),
   277 => (x"da",x"c1",x"87",x"df"),
   278 => (x"87",x"fd",x"e1",x"49"),
   279 => (x"f8",x"c2",x"4d",x"c1"),
   280 => (x"02",x"bf",x"97",x"c4"),
   281 => (x"db",x"c2",x"87",x"cf"),
   282 => (x"c1",x"49",x"bf",x"da"),
   283 => (x"de",x"db",x"c2",x"b9"),
   284 => (x"cf",x"fa",x"71",x"59"),
   285 => (x"c9",x"f8",x"c2",x"87"),
   286 => (x"db",x"c2",x"4b",x"bf"),
   287 => (x"c1",x"05",x"bf",x"f6"),
   288 => (x"db",x"c2",x"87",x"e1"),
   289 => (x"c0",x"02",x"bf",x"de"),
   290 => (x"a6",x"c4",x"87",x"f0"),
   291 => (x"c0",x"c0",x"c8",x"48"),
   292 => (x"e2",x"db",x"c2",x"78"),
   293 => (x"bf",x"97",x"6e",x"7e"),
   294 => (x"c1",x"48",x"6e",x"49"),
   295 => (x"71",x"7e",x"70",x"80"),
   296 => (x"70",x"87",x"f6",x"e0"),
   297 => (x"87",x"c3",x"02",x"98"),
   298 => (x"c4",x"b3",x"66",x"c4"),
   299 => (x"b7",x"c1",x"48",x"66"),
   300 => (x"58",x"a6",x"c8",x"28"),
   301 => (x"ff",x"05",x"98",x"70"),
   302 => (x"fd",x"c3",x"87",x"db"),
   303 => (x"87",x"d9",x"e0",x"49"),
   304 => (x"e0",x"49",x"fa",x"c3"),
   305 => (x"49",x"73",x"87",x"d3"),
   306 => (x"71",x"99",x"ff",x"c3"),
   307 => (x"f8",x"49",x"c0",x"1e"),
   308 => (x"49",x"73",x"87",x"e4"),
   309 => (x"71",x"29",x"b7",x"c8"),
   310 => (x"f8",x"49",x"c1",x"1e"),
   311 => (x"86",x"c8",x"87",x"d8"),
   312 => (x"c2",x"87",x"c9",x"c6"),
   313 => (x"4b",x"bf",x"cd",x"f8"),
   314 => (x"87",x"df",x"02",x"9b"),
   315 => (x"bf",x"f2",x"db",x"c2"),
   316 => (x"87",x"d6",x"c8",x"49"),
   317 => (x"c0",x"05",x"98",x"70"),
   318 => (x"4b",x"c0",x"87",x"c4"),
   319 => (x"e0",x"c2",x"87",x"d3"),
   320 => (x"87",x"fa",x"c7",x"49"),
   321 => (x"58",x"f6",x"db",x"c2"),
   322 => (x"c2",x"87",x"c6",x"c0"),
   323 => (x"c0",x"48",x"f2",x"db"),
   324 => (x"c2",x"49",x"73",x"78"),
   325 => (x"cf",x"c0",x"05",x"99"),
   326 => (x"49",x"eb",x"c3",x"87"),
   327 => (x"87",x"f9",x"de",x"ff"),
   328 => (x"99",x"c2",x"49",x"70"),
   329 => (x"87",x"c2",x"c0",x"02"),
   330 => (x"49",x"73",x"4c",x"fb"),
   331 => (x"c0",x"05",x"99",x"c1"),
   332 => (x"f4",x"c3",x"87",x"cf"),
   333 => (x"e0",x"de",x"ff",x"49"),
   334 => (x"c2",x"49",x"70",x"87"),
   335 => (x"c2",x"c0",x"02",x"99"),
   336 => (x"73",x"4c",x"fa",x"87"),
   337 => (x"05",x"99",x"c8",x"49"),
   338 => (x"c3",x"87",x"cf",x"c0"),
   339 => (x"de",x"ff",x"49",x"f5"),
   340 => (x"49",x"70",x"87",x"c7"),
   341 => (x"c0",x"02",x"99",x"c2"),
   342 => (x"f8",x"c2",x"87",x"d6"),
   343 => (x"c0",x"02",x"bf",x"d5"),
   344 => (x"c1",x"48",x"87",x"ca"),
   345 => (x"d9",x"f8",x"c2",x"88"),
   346 => (x"87",x"c2",x"c0",x"58"),
   347 => (x"4d",x"c1",x"4c",x"ff"),
   348 => (x"99",x"c4",x"49",x"73"),
   349 => (x"87",x"cf",x"c0",x"05"),
   350 => (x"ff",x"49",x"f2",x"c3"),
   351 => (x"70",x"87",x"da",x"dd"),
   352 => (x"02",x"99",x"c2",x"49"),
   353 => (x"c2",x"87",x"dc",x"c0"),
   354 => (x"7e",x"bf",x"d5",x"f8"),
   355 => (x"a8",x"b7",x"c7",x"48"),
   356 => (x"87",x"cb",x"c0",x"03"),
   357 => (x"80",x"c1",x"48",x"6e"),
   358 => (x"58",x"d9",x"f8",x"c2"),
   359 => (x"fe",x"87",x"c2",x"c0"),
   360 => (x"c3",x"4d",x"c1",x"4c"),
   361 => (x"dc",x"ff",x"49",x"fd"),
   362 => (x"49",x"70",x"87",x"ef"),
   363 => (x"c0",x"02",x"99",x"c2"),
   364 => (x"f8",x"c2",x"87",x"d5"),
   365 => (x"c0",x"02",x"bf",x"d5"),
   366 => (x"f8",x"c2",x"87",x"c9"),
   367 => (x"78",x"c0",x"48",x"d5"),
   368 => (x"fd",x"87",x"c2",x"c0"),
   369 => (x"c3",x"4d",x"c1",x"4c"),
   370 => (x"dc",x"ff",x"49",x"fa"),
   371 => (x"49",x"70",x"87",x"cb"),
   372 => (x"c0",x"02",x"99",x"c2"),
   373 => (x"f8",x"c2",x"87",x"d9"),
   374 => (x"c7",x"48",x"bf",x"d5"),
   375 => (x"c0",x"03",x"a8",x"b7"),
   376 => (x"f8",x"c2",x"87",x"c9"),
   377 => (x"78",x"c7",x"48",x"d5"),
   378 => (x"fc",x"87",x"c2",x"c0"),
   379 => (x"c0",x"4d",x"c1",x"4c"),
   380 => (x"c0",x"03",x"ac",x"b7"),
   381 => (x"66",x"c4",x"87",x"d0"),
   382 => (x"82",x"d8",x"c1",x"4a"),
   383 => (x"c5",x"c0",x"02",x"6a"),
   384 => (x"49",x"74",x"4b",x"87"),
   385 => (x"1e",x"c0",x"0f",x"73"),
   386 => (x"c1",x"1e",x"f0",x"c3"),
   387 => (x"c2",x"f5",x"49",x"da"),
   388 => (x"70",x"86",x"c8",x"87"),
   389 => (x"e0",x"c0",x"02",x"98"),
   390 => (x"48",x"a6",x"c8",x"87"),
   391 => (x"bf",x"d5",x"f8",x"c2"),
   392 => (x"49",x"66",x"c8",x"78"),
   393 => (x"66",x"c4",x"91",x"cb"),
   394 => (x"70",x"80",x"71",x"48"),
   395 => (x"02",x"bf",x"6e",x"7e"),
   396 => (x"4b",x"87",x"c6",x"c0"),
   397 => (x"73",x"49",x"66",x"c8"),
   398 => (x"02",x"9d",x"75",x"0f"),
   399 => (x"c2",x"87",x"c8",x"c0"),
   400 => (x"49",x"bf",x"d5",x"f8"),
   401 => (x"c2",x"87",x"c9",x"f0"),
   402 => (x"02",x"bf",x"fa",x"db"),
   403 => (x"49",x"87",x"dd",x"c0"),
   404 => (x"70",x"87",x"f7",x"c2"),
   405 => (x"d3",x"c0",x"02",x"98"),
   406 => (x"d5",x"f8",x"c2",x"87"),
   407 => (x"ef",x"ef",x"49",x"bf"),
   408 => (x"f1",x"49",x"c0",x"87"),
   409 => (x"db",x"c2",x"87",x"cf"),
   410 => (x"78",x"c0",x"48",x"fa"),
   411 => (x"e9",x"f0",x"8e",x"f4"),
   412 => (x"79",x"6f",x"4a",x"87"),
   413 => (x"73",x"79",x"65",x"6b"),
   414 => (x"00",x"6e",x"6f",x"20"),
   415 => (x"6b",x"79",x"6f",x"4a"),
   416 => (x"20",x"73",x"79",x"65"),
   417 => (x"00",x"66",x"66",x"6f"),
   418 => (x"5c",x"5b",x"5e",x"0e"),
   419 => (x"71",x"1e",x"0e",x"5d"),
   420 => (x"d1",x"f8",x"c2",x"4c"),
   421 => (x"cd",x"c1",x"49",x"bf"),
   422 => (x"d1",x"c1",x"4d",x"a1"),
   423 => (x"74",x"7e",x"69",x"81"),
   424 => (x"87",x"cf",x"02",x"9c"),
   425 => (x"74",x"4b",x"a5",x"c4"),
   426 => (x"d1",x"f8",x"c2",x"7b"),
   427 => (x"f1",x"ef",x"49",x"bf"),
   428 => (x"74",x"7b",x"6e",x"87"),
   429 => (x"87",x"c4",x"05",x"9c"),
   430 => (x"87",x"c2",x"4b",x"c0"),
   431 => (x"49",x"73",x"4b",x"c1"),
   432 => (x"d4",x"87",x"f2",x"ef"),
   433 => (x"87",x"c8",x"02",x"66"),
   434 => (x"87",x"f2",x"c0",x"49"),
   435 => (x"87",x"c2",x"4a",x"70"),
   436 => (x"db",x"c2",x"4a",x"c0"),
   437 => (x"ef",x"26",x"5a",x"fe"),
   438 => (x"00",x"00",x"87",x"c0"),
   439 => (x"00",x"00",x"00",x"00"),
   440 => (x"12",x"58",x"00",x"00"),
   441 => (x"1b",x"1d",x"14",x"11"),
   442 => (x"59",x"5a",x"23",x"1c"),
   443 => (x"f2",x"f5",x"94",x"91"),
   444 => (x"00",x"00",x"f4",x"eb"),
   445 => (x"00",x"00",x"00",x"00"),
   446 => (x"00",x"00",x"00",x"00"),
   447 => (x"71",x"1e",x"00",x"00"),
   448 => (x"bf",x"c8",x"ff",x"4a"),
   449 => (x"48",x"a1",x"72",x"49"),
   450 => (x"ff",x"1e",x"4f",x"26"),
   451 => (x"fe",x"89",x"bf",x"c8"),
   452 => (x"c0",x"c0",x"c0",x"c0"),
   453 => (x"c4",x"01",x"a9",x"c0"),
   454 => (x"c2",x"4a",x"c0",x"87"),
   455 => (x"72",x"4a",x"c1",x"87"),
   456 => (x"0e",x"4f",x"26",x"48"),
   457 => (x"5d",x"5c",x"5b",x"5e"),
   458 => (x"ff",x"4b",x"71",x"0e"),
   459 => (x"66",x"d0",x"4c",x"d4"),
   460 => (x"d6",x"78",x"c0",x"48"),
   461 => (x"d8",x"d8",x"ff",x"49"),
   462 => (x"7c",x"ff",x"c3",x"87"),
   463 => (x"ff",x"c3",x"49",x"6c"),
   464 => (x"49",x"4d",x"71",x"99"),
   465 => (x"c1",x"99",x"f0",x"c3"),
   466 => (x"cb",x"05",x"a9",x"e0"),
   467 => (x"7c",x"ff",x"c3",x"87"),
   468 => (x"98",x"c3",x"48",x"6c"),
   469 => (x"78",x"08",x"66",x"d0"),
   470 => (x"6c",x"7c",x"ff",x"c3"),
   471 => (x"31",x"c8",x"49",x"4a"),
   472 => (x"6c",x"7c",x"ff",x"c3"),
   473 => (x"72",x"b2",x"71",x"4a"),
   474 => (x"c3",x"31",x"c8",x"49"),
   475 => (x"4a",x"6c",x"7c",x"ff"),
   476 => (x"49",x"72",x"b2",x"71"),
   477 => (x"ff",x"c3",x"31",x"c8"),
   478 => (x"71",x"4a",x"6c",x"7c"),
   479 => (x"48",x"d0",x"ff",x"b2"),
   480 => (x"73",x"78",x"e0",x"c0"),
   481 => (x"87",x"c2",x"02",x"9b"),
   482 => (x"48",x"75",x"7b",x"72"),
   483 => (x"4c",x"26",x"4d",x"26"),
   484 => (x"4f",x"26",x"4b",x"26"),
   485 => (x"0e",x"4f",x"26",x"1e"),
   486 => (x"0e",x"5c",x"5b",x"5e"),
   487 => (x"1e",x"76",x"86",x"f8"),
   488 => (x"fd",x"49",x"a6",x"c8"),
   489 => (x"86",x"c4",x"87",x"fd"),
   490 => (x"48",x"6e",x"4b",x"70"),
   491 => (x"c2",x"03",x"a8",x"c2"),
   492 => (x"4a",x"73",x"87",x"f0"),
   493 => (x"c1",x"9a",x"f0",x"c3"),
   494 => (x"c7",x"02",x"aa",x"d0"),
   495 => (x"aa",x"e0",x"c1",x"87"),
   496 => (x"87",x"de",x"c2",x"05"),
   497 => (x"99",x"c8",x"49",x"73"),
   498 => (x"ff",x"87",x"c3",x"02"),
   499 => (x"4c",x"73",x"87",x"c6"),
   500 => (x"ac",x"c2",x"9c",x"c3"),
   501 => (x"87",x"c2",x"c1",x"05"),
   502 => (x"c9",x"49",x"66",x"c4"),
   503 => (x"c4",x"1e",x"71",x"31"),
   504 => (x"92",x"d4",x"4a",x"66"),
   505 => (x"49",x"d9",x"f8",x"c2"),
   506 => (x"c7",x"fe",x"81",x"72"),
   507 => (x"49",x"d8",x"87",x"e4"),
   508 => (x"87",x"dd",x"d5",x"ff"),
   509 => (x"c2",x"1e",x"c0",x"c8"),
   510 => (x"fd",x"49",x"f6",x"e6"),
   511 => (x"ff",x"87",x"df",x"e3"),
   512 => (x"e0",x"c0",x"48",x"d0"),
   513 => (x"f6",x"e6",x"c2",x"78"),
   514 => (x"4a",x"66",x"cc",x"1e"),
   515 => (x"f8",x"c2",x"92",x"d4"),
   516 => (x"81",x"72",x"49",x"d9"),
   517 => (x"87",x"eb",x"c5",x"fe"),
   518 => (x"ac",x"c1",x"86",x"cc"),
   519 => (x"87",x"c2",x"c1",x"05"),
   520 => (x"c9",x"49",x"66",x"c4"),
   521 => (x"c4",x"1e",x"71",x"31"),
   522 => (x"92",x"d4",x"4a",x"66"),
   523 => (x"49",x"d9",x"f8",x"c2"),
   524 => (x"c6",x"fe",x"81",x"72"),
   525 => (x"e6",x"c2",x"87",x"dc"),
   526 => (x"66",x"c8",x"1e",x"f6"),
   527 => (x"c2",x"92",x"d4",x"4a"),
   528 => (x"72",x"49",x"d9",x"f8"),
   529 => (x"eb",x"c3",x"fe",x"81"),
   530 => (x"ff",x"49",x"d7",x"87"),
   531 => (x"c8",x"87",x"c2",x"d4"),
   532 => (x"e6",x"c2",x"1e",x"c0"),
   533 => (x"e1",x"fd",x"49",x"f6"),
   534 => (x"86",x"cc",x"87",x"dd"),
   535 => (x"c0",x"48",x"d0",x"ff"),
   536 => (x"8e",x"f8",x"78",x"e0"),
   537 => (x"0e",x"87",x"e7",x"fc"),
   538 => (x"5d",x"5c",x"5b",x"5e"),
   539 => (x"4d",x"71",x"1e",x"0e"),
   540 => (x"d4",x"4c",x"d4",x"ff"),
   541 => (x"c3",x"48",x"7e",x"66"),
   542 => (x"c5",x"06",x"a8",x"b7"),
   543 => (x"c1",x"48",x"c0",x"87"),
   544 => (x"49",x"75",x"87",x"e2"),
   545 => (x"87",x"d7",x"d4",x"fe"),
   546 => (x"66",x"c4",x"1e",x"75"),
   547 => (x"c2",x"93",x"d4",x"4b"),
   548 => (x"73",x"83",x"d9",x"f8"),
   549 => (x"e7",x"fd",x"fd",x"49"),
   550 => (x"6b",x"83",x"c8",x"87"),
   551 => (x"48",x"d0",x"ff",x"4b"),
   552 => (x"dd",x"78",x"e1",x"c8"),
   553 => (x"c3",x"49",x"73",x"7c"),
   554 => (x"7c",x"71",x"99",x"ff"),
   555 => (x"b7",x"c8",x"49",x"73"),
   556 => (x"99",x"ff",x"c3",x"29"),
   557 => (x"49",x"73",x"7c",x"71"),
   558 => (x"c3",x"29",x"b7",x"d0"),
   559 => (x"7c",x"71",x"99",x"ff"),
   560 => (x"b7",x"d8",x"49",x"73"),
   561 => (x"c0",x"7c",x"71",x"29"),
   562 => (x"7c",x"7c",x"7c",x"7c"),
   563 => (x"7c",x"7c",x"7c",x"7c"),
   564 => (x"7c",x"7c",x"7c",x"7c"),
   565 => (x"c4",x"78",x"e0",x"c0"),
   566 => (x"49",x"dc",x"1e",x"66"),
   567 => (x"87",x"d6",x"d2",x"ff"),
   568 => (x"48",x"73",x"86",x"c8"),
   569 => (x"87",x"e4",x"fa",x"26"),
   570 => (x"c4",x"4a",x"71",x"1e"),
   571 => (x"f7",x"c2",x"49",x"a2"),
   572 => (x"78",x"6a",x"48",x"f0"),
   573 => (x"48",x"da",x"db",x"c2"),
   574 => (x"db",x"c2",x"78",x"69"),
   575 => (x"e8",x"49",x"bf",x"da"),
   576 => (x"d3",x"ff",x"87",x"c2"),
   577 => (x"48",x"c1",x"87",x"ca"),
   578 => (x"71",x"1e",x"4f",x"26"),
   579 => (x"49",x"a2",x"c4",x"4a"),
   580 => (x"bf",x"f0",x"f7",x"c2"),
   581 => (x"da",x"db",x"c2",x"7a"),
   582 => (x"4f",x"26",x"79",x"bf"),
   583 => (x"9a",x"4a",x"71",x"1e"),
   584 => (x"87",x"ec",x"c0",x"02"),
   585 => (x"ec",x"f3",x"c2",x"1e"),
   586 => (x"d3",x"fb",x"fd",x"49"),
   587 => (x"70",x"86",x"c4",x"87"),
   588 => (x"87",x"dc",x"02",x"98"),
   589 => (x"1e",x"f6",x"e6",x"c2"),
   590 => (x"49",x"ec",x"f3",x"c2"),
   591 => (x"87",x"f4",x"ff",x"fd"),
   592 => (x"98",x"70",x"86",x"c4"),
   593 => (x"c2",x"87",x"c9",x"02"),
   594 => (x"fe",x"49",x"f6",x"e6"),
   595 => (x"87",x"c2",x"87",x"da"),
   596 => (x"4f",x"26",x"48",x"c0"),
   597 => (x"9a",x"4a",x"71",x"1e"),
   598 => (x"87",x"ee",x"c0",x"02"),
   599 => (x"ec",x"f3",x"c2",x"1e"),
   600 => (x"db",x"fa",x"fd",x"49"),
   601 => (x"70",x"86",x"c4",x"87"),
   602 => (x"87",x"de",x"02",x"98"),
   603 => (x"49",x"f6",x"e6",x"c2"),
   604 => (x"c2",x"87",x"d7",x"fe"),
   605 => (x"c2",x"1e",x"f6",x"e6"),
   606 => (x"fe",x"49",x"ec",x"f3"),
   607 => (x"c4",x"87",x"c4",x"c0"),
   608 => (x"02",x"98",x"70",x"86"),
   609 => (x"48",x"c1",x"87",x"c4"),
   610 => (x"48",x"c0",x"87",x"c2"),
   611 => (x"48",x"c0",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

