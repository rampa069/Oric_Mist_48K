
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"ff",x"cf",x"87",x"c4"),
     1 => (x"fb",x"c2",x"4a",x"ff"),
     2 => (x"fb",x"c2",x"5a",x"c0"),
     3 => (x"78",x"c1",x"48",x"c0"),
     4 => (x"4f",x"26",x"4b",x"26"),
     5 => (x"5c",x"5b",x"5e",x"0e"),
     6 => (x"4d",x"71",x"0e",x"5d"),
     7 => (x"bf",x"fc",x"fa",x"c2"),
     8 => (x"02",x"9d",x"75",x"4b"),
     9 => (x"c8",x"49",x"87",x"cb"),
    10 => (x"fc",x"fe",x"c1",x"91"),
    11 => (x"c4",x"82",x"71",x"4a"),
    12 => (x"fc",x"c2",x"c2",x"87"),
    13 => (x"12",x"4c",x"c0",x"4a"),
    14 => (x"c2",x"99",x"73",x"49"),
    15 => (x"48",x"bf",x"f8",x"fa"),
    16 => (x"d4",x"ff",x"b8",x"71"),
    17 => (x"b7",x"c1",x"78",x"08"),
    18 => (x"b7",x"c8",x"84",x"2b"),
    19 => (x"87",x"e7",x"04",x"ac"),
    20 => (x"bf",x"f4",x"fa",x"c2"),
    21 => (x"c2",x"80",x"c8",x"48"),
    22 => (x"26",x"58",x"f8",x"fa"),
    23 => (x"26",x"4c",x"26",x"4d"),
    24 => (x"1e",x"4f",x"26",x"4b"),
    25 => (x"4b",x"71",x"1e",x"73"),
    26 => (x"02",x"9a",x"4a",x"13"),
    27 => (x"49",x"72",x"87",x"cb"),
    28 => (x"13",x"87",x"e1",x"fe"),
    29 => (x"f5",x"05",x"9a",x"4a"),
    30 => (x"26",x"4b",x"26",x"87"),
    31 => (x"fa",x"c2",x"1e",x"4f"),
    32 => (x"c2",x"49",x"bf",x"f4"),
    33 => (x"c1",x"48",x"f4",x"fa"),
    34 => (x"c0",x"c4",x"78",x"a1"),
    35 => (x"db",x"03",x"a9",x"b7"),
    36 => (x"48",x"d4",x"ff",x"87"),
    37 => (x"bf",x"f8",x"fa",x"c2"),
    38 => (x"f4",x"fa",x"c2",x"78"),
    39 => (x"fa",x"c2",x"49",x"bf"),
    40 => (x"a1",x"c1",x"48",x"f4"),
    41 => (x"b7",x"c0",x"c4",x"78"),
    42 => (x"87",x"e5",x"04",x"a9"),
    43 => (x"c8",x"48",x"d0",x"ff"),
    44 => (x"c0",x"fb",x"c2",x"78"),
    45 => (x"26",x"78",x"c0",x"48"),
    46 => (x"00",x"00",x"00",x"4f"),
    47 => (x"00",x"00",x"00",x"00"),
    48 => (x"00",x"00",x"00",x"00"),
    49 => (x"5f",x"00",x"00",x"00"),
    50 => (x"00",x"00",x"00",x"5f"),
    51 => (x"00",x"03",x"03",x"00"),
    52 => (x"00",x"00",x"03",x"03"),
    53 => (x"14",x"7f",x"7f",x"14"),
    54 => (x"00",x"14",x"7f",x"7f"),
    55 => (x"6b",x"2e",x"24",x"00"),
    56 => (x"00",x"12",x"3a",x"6b"),
    57 => (x"18",x"36",x"6a",x"4c"),
    58 => (x"00",x"32",x"56",x"6c"),
    59 => (x"59",x"4f",x"7e",x"30"),
    60 => (x"40",x"68",x"3a",x"77"),
    61 => (x"07",x"04",x"00",x"00"),
    62 => (x"00",x"00",x"00",x"03"),
    63 => (x"3e",x"1c",x"00",x"00"),
    64 => (x"00",x"00",x"41",x"63"),
    65 => (x"63",x"41",x"00",x"00"),
    66 => (x"00",x"00",x"1c",x"3e"),
    67 => (x"1c",x"3e",x"2a",x"08"),
    68 => (x"08",x"2a",x"3e",x"1c"),
    69 => (x"3e",x"08",x"08",x"00"),
    70 => (x"00",x"08",x"08",x"3e"),
    71 => (x"e0",x"80",x"00",x"00"),
    72 => (x"00",x"00",x"00",x"60"),
    73 => (x"08",x"08",x"08",x"00"),
    74 => (x"00",x"08",x"08",x"08"),
    75 => (x"60",x"00",x"00",x"00"),
    76 => (x"00",x"00",x"00",x"60"),
    77 => (x"18",x"30",x"60",x"40"),
    78 => (x"01",x"03",x"06",x"0c"),
    79 => (x"59",x"7f",x"3e",x"00"),
    80 => (x"00",x"3e",x"7f",x"4d"),
    81 => (x"7f",x"06",x"04",x"00"),
    82 => (x"00",x"00",x"00",x"7f"),
    83 => (x"71",x"63",x"42",x"00"),
    84 => (x"00",x"46",x"4f",x"59"),
    85 => (x"49",x"63",x"22",x"00"),
    86 => (x"00",x"36",x"7f",x"49"),
    87 => (x"13",x"16",x"1c",x"18"),
    88 => (x"00",x"10",x"7f",x"7f"),
    89 => (x"45",x"67",x"27",x"00"),
    90 => (x"00",x"39",x"7d",x"45"),
    91 => (x"4b",x"7e",x"3c",x"00"),
    92 => (x"00",x"30",x"79",x"49"),
    93 => (x"71",x"01",x"01",x"00"),
    94 => (x"00",x"07",x"0f",x"79"),
    95 => (x"49",x"7f",x"36",x"00"),
    96 => (x"00",x"36",x"7f",x"49"),
    97 => (x"49",x"4f",x"06",x"00"),
    98 => (x"00",x"1e",x"3f",x"69"),
    99 => (x"66",x"00",x"00",x"00"),
   100 => (x"00",x"00",x"00",x"66"),
   101 => (x"e6",x"80",x"00",x"00"),
   102 => (x"00",x"00",x"00",x"66"),
   103 => (x"14",x"08",x"08",x"00"),
   104 => (x"00",x"22",x"22",x"14"),
   105 => (x"14",x"14",x"14",x"00"),
   106 => (x"00",x"14",x"14",x"14"),
   107 => (x"14",x"22",x"22",x"00"),
   108 => (x"00",x"08",x"08",x"14"),
   109 => (x"51",x"03",x"02",x"00"),
   110 => (x"00",x"06",x"0f",x"59"),
   111 => (x"5d",x"41",x"7f",x"3e"),
   112 => (x"00",x"1e",x"1f",x"55"),
   113 => (x"09",x"7f",x"7e",x"00"),
   114 => (x"00",x"7e",x"7f",x"09"),
   115 => (x"49",x"7f",x"7f",x"00"),
   116 => (x"00",x"36",x"7f",x"49"),
   117 => (x"63",x"3e",x"1c",x"00"),
   118 => (x"00",x"41",x"41",x"41"),
   119 => (x"41",x"7f",x"7f",x"00"),
   120 => (x"00",x"1c",x"3e",x"63"),
   121 => (x"49",x"7f",x"7f",x"00"),
   122 => (x"00",x"41",x"41",x"49"),
   123 => (x"09",x"7f",x"7f",x"00"),
   124 => (x"00",x"01",x"01",x"09"),
   125 => (x"41",x"7f",x"3e",x"00"),
   126 => (x"00",x"7a",x"7b",x"49"),
   127 => (x"08",x"7f",x"7f",x"00"),
   128 => (x"00",x"7f",x"7f",x"08"),
   129 => (x"7f",x"41",x"00",x"00"),
   130 => (x"00",x"00",x"41",x"7f"),
   131 => (x"40",x"60",x"20",x"00"),
   132 => (x"00",x"3f",x"7f",x"40"),
   133 => (x"1c",x"08",x"7f",x"7f"),
   134 => (x"00",x"41",x"63",x"36"),
   135 => (x"40",x"7f",x"7f",x"00"),
   136 => (x"00",x"40",x"40",x"40"),
   137 => (x"0c",x"06",x"7f",x"7f"),
   138 => (x"00",x"7f",x"7f",x"06"),
   139 => (x"0c",x"06",x"7f",x"7f"),
   140 => (x"00",x"7f",x"7f",x"18"),
   141 => (x"41",x"7f",x"3e",x"00"),
   142 => (x"00",x"3e",x"7f",x"41"),
   143 => (x"09",x"7f",x"7f",x"00"),
   144 => (x"00",x"06",x"0f",x"09"),
   145 => (x"61",x"41",x"7f",x"3e"),
   146 => (x"00",x"40",x"7e",x"7f"),
   147 => (x"09",x"7f",x"7f",x"00"),
   148 => (x"00",x"66",x"7f",x"19"),
   149 => (x"4d",x"6f",x"26",x"00"),
   150 => (x"00",x"32",x"7b",x"59"),
   151 => (x"7f",x"01",x"01",x"00"),
   152 => (x"00",x"01",x"01",x"7f"),
   153 => (x"40",x"7f",x"3f",x"00"),
   154 => (x"00",x"3f",x"7f",x"40"),
   155 => (x"70",x"3f",x"0f",x"00"),
   156 => (x"00",x"0f",x"3f",x"70"),
   157 => (x"18",x"30",x"7f",x"7f"),
   158 => (x"00",x"7f",x"7f",x"30"),
   159 => (x"1c",x"36",x"63",x"41"),
   160 => (x"41",x"63",x"36",x"1c"),
   161 => (x"7c",x"06",x"03",x"01"),
   162 => (x"01",x"03",x"06",x"7c"),
   163 => (x"4d",x"59",x"71",x"61"),
   164 => (x"00",x"41",x"43",x"47"),
   165 => (x"7f",x"7f",x"00",x"00"),
   166 => (x"00",x"00",x"41",x"41"),
   167 => (x"0c",x"06",x"03",x"01"),
   168 => (x"40",x"60",x"30",x"18"),
   169 => (x"41",x"41",x"00",x"00"),
   170 => (x"00",x"00",x"7f",x"7f"),
   171 => (x"03",x"06",x"0c",x"08"),
   172 => (x"00",x"08",x"0c",x"06"),
   173 => (x"80",x"80",x"80",x"80"),
   174 => (x"00",x"80",x"80",x"80"),
   175 => (x"03",x"00",x"00",x"00"),
   176 => (x"00",x"00",x"04",x"07"),
   177 => (x"54",x"74",x"20",x"00"),
   178 => (x"00",x"78",x"7c",x"54"),
   179 => (x"44",x"7f",x"7f",x"00"),
   180 => (x"00",x"38",x"7c",x"44"),
   181 => (x"44",x"7c",x"38",x"00"),
   182 => (x"00",x"00",x"44",x"44"),
   183 => (x"44",x"7c",x"38",x"00"),
   184 => (x"00",x"7f",x"7f",x"44"),
   185 => (x"54",x"7c",x"38",x"00"),
   186 => (x"00",x"18",x"5c",x"54"),
   187 => (x"7f",x"7e",x"04",x"00"),
   188 => (x"00",x"00",x"05",x"05"),
   189 => (x"a4",x"bc",x"18",x"00"),
   190 => (x"00",x"7c",x"fc",x"a4"),
   191 => (x"04",x"7f",x"7f",x"00"),
   192 => (x"00",x"78",x"7c",x"04"),
   193 => (x"3d",x"00",x"00",x"00"),
   194 => (x"00",x"00",x"40",x"7d"),
   195 => (x"80",x"80",x"80",x"00"),
   196 => (x"00",x"00",x"7d",x"fd"),
   197 => (x"10",x"7f",x"7f",x"00"),
   198 => (x"00",x"44",x"6c",x"38"),
   199 => (x"3f",x"00",x"00",x"00"),
   200 => (x"00",x"00",x"40",x"7f"),
   201 => (x"18",x"0c",x"7c",x"7c"),
   202 => (x"00",x"78",x"7c",x"0c"),
   203 => (x"04",x"7c",x"7c",x"00"),
   204 => (x"00",x"78",x"7c",x"04"),
   205 => (x"44",x"7c",x"38",x"00"),
   206 => (x"00",x"38",x"7c",x"44"),
   207 => (x"24",x"fc",x"fc",x"00"),
   208 => (x"00",x"18",x"3c",x"24"),
   209 => (x"24",x"3c",x"18",x"00"),
   210 => (x"00",x"fc",x"fc",x"24"),
   211 => (x"04",x"7c",x"7c",x"00"),
   212 => (x"00",x"08",x"0c",x"04"),
   213 => (x"54",x"5c",x"48",x"00"),
   214 => (x"00",x"20",x"74",x"54"),
   215 => (x"7f",x"3f",x"04",x"00"),
   216 => (x"00",x"00",x"44",x"44"),
   217 => (x"40",x"7c",x"3c",x"00"),
   218 => (x"00",x"7c",x"7c",x"40"),
   219 => (x"60",x"3c",x"1c",x"00"),
   220 => (x"00",x"1c",x"3c",x"60"),
   221 => (x"30",x"60",x"7c",x"3c"),
   222 => (x"00",x"3c",x"7c",x"60"),
   223 => (x"10",x"38",x"6c",x"44"),
   224 => (x"00",x"44",x"6c",x"38"),
   225 => (x"e0",x"bc",x"1c",x"00"),
   226 => (x"00",x"1c",x"3c",x"60"),
   227 => (x"74",x"64",x"44",x"00"),
   228 => (x"00",x"44",x"4c",x"5c"),
   229 => (x"3e",x"08",x"08",x"00"),
   230 => (x"00",x"41",x"41",x"77"),
   231 => (x"7f",x"00",x"00",x"00"),
   232 => (x"00",x"00",x"00",x"7f"),
   233 => (x"77",x"41",x"41",x"00"),
   234 => (x"00",x"08",x"08",x"3e"),
   235 => (x"03",x"01",x"01",x"02"),
   236 => (x"00",x"01",x"02",x"02"),
   237 => (x"7f",x"7f",x"7f",x"7f"),
   238 => (x"00",x"7f",x"7f",x"7f"),
   239 => (x"1c",x"1c",x"08",x"08"),
   240 => (x"7f",x"7f",x"3e",x"3e"),
   241 => (x"3e",x"3e",x"7f",x"7f"),
   242 => (x"08",x"08",x"1c",x"1c"),
   243 => (x"7c",x"18",x"10",x"00"),
   244 => (x"00",x"10",x"18",x"7c"),
   245 => (x"7c",x"30",x"10",x"00"),
   246 => (x"00",x"10",x"30",x"7c"),
   247 => (x"60",x"60",x"30",x"10"),
   248 => (x"00",x"06",x"1e",x"78"),
   249 => (x"18",x"3c",x"66",x"42"),
   250 => (x"00",x"42",x"66",x"3c"),
   251 => (x"c2",x"6a",x"38",x"78"),
   252 => (x"00",x"38",x"6c",x"c6"),
   253 => (x"60",x"00",x"00",x"60"),
   254 => (x"00",x"60",x"00",x"00"),
   255 => (x"5c",x"5b",x"5e",x"0e"),
   256 => (x"86",x"fc",x"0e",x"5d"),
   257 => (x"fb",x"c2",x"7e",x"71"),
   258 => (x"c0",x"4c",x"bf",x"c8"),
   259 => (x"c4",x"1e",x"c0",x"4b"),
   260 => (x"c4",x"02",x"ab",x"66"),
   261 => (x"c2",x"4d",x"c0",x"87"),
   262 => (x"75",x"4d",x"c1",x"87"),
   263 => (x"ee",x"49",x"73",x"1e"),
   264 => (x"86",x"c8",x"87",x"e1"),
   265 => (x"ef",x"49",x"e0",x"c0"),
   266 => (x"a4",x"c4",x"87",x"ea"),
   267 => (x"f0",x"49",x"6a",x"4a"),
   268 => (x"c8",x"f1",x"87",x"f1"),
   269 => (x"c1",x"84",x"cc",x"87"),
   270 => (x"ab",x"b7",x"c8",x"83"),
   271 => (x"87",x"cd",x"ff",x"04"),
   272 => (x"4d",x"26",x"8e",x"fc"),
   273 => (x"4b",x"26",x"4c",x"26"),
   274 => (x"71",x"1e",x"4f",x"26"),
   275 => (x"cc",x"fb",x"c2",x"4a"),
   276 => (x"cc",x"fb",x"c2",x"5a"),
   277 => (x"49",x"78",x"c7",x"48"),
   278 => (x"26",x"87",x"e1",x"fe"),
   279 => (x"1e",x"73",x"1e",x"4f"),
   280 => (x"0b",x"fc",x"4b",x"71"),
   281 => (x"4a",x"73",x"0b",x"7b"),
   282 => (x"c0",x"c1",x"9a",x"c1"),
   283 => (x"c5",x"ed",x"49",x"a2"),
   284 => (x"cc",x"df",x"c2",x"87"),
   285 => (x"26",x"4b",x"26",x"5b"),
   286 => (x"4a",x"71",x"1e",x"4f"),
   287 => (x"72",x"1e",x"66",x"c4"),
   288 => (x"87",x"cb",x"ec",x"49"),
   289 => (x"4f",x"26",x"8e",x"fc"),
   290 => (x"48",x"d4",x"ff",x"1e"),
   291 => (x"ff",x"78",x"ff",x"c3"),
   292 => (x"e1",x"c0",x"48",x"d0"),
   293 => (x"48",x"d4",x"ff",x"78"),
   294 => (x"48",x"71",x"78",x"c1"),
   295 => (x"d4",x"ff",x"30",x"c4"),
   296 => (x"d0",x"ff",x"78",x"08"),
   297 => (x"78",x"e0",x"c0",x"48"),
   298 => (x"5e",x"0e",x"4f",x"26"),
   299 => (x"0e",x"5d",x"5c",x"5b"),
   300 => (x"a6",x"c8",x"86",x"ec"),
   301 => (x"c4",x"78",x"c0",x"48"),
   302 => (x"78",x"bf",x"ec",x"80"),
   303 => (x"fb",x"c2",x"80",x"f8"),
   304 => (x"c2",x"78",x"bf",x"c8"),
   305 => (x"4c",x"bf",x"d0",x"fb"),
   306 => (x"c2",x"4d",x"bf",x"e8"),
   307 => (x"49",x"bf",x"c8",x"df"),
   308 => (x"c7",x"87",x"c7",x"e4"),
   309 => (x"87",x"ff",x"e8",x"49"),
   310 => (x"99",x"c2",x"49",x"70"),
   311 => (x"c2",x"87",x"d0",x"05"),
   312 => (x"49",x"bf",x"c0",x"df"),
   313 => (x"66",x"cc",x"b9",x"ff"),
   314 => (x"02",x"99",x"c1",x"99"),
   315 => (x"c8",x"87",x"cb",x"c2"),
   316 => (x"c8",x"ff",x"48",x"a6"),
   317 => (x"49",x"c7",x"78",x"bf"),
   318 => (x"70",x"87",x"dc",x"e8"),
   319 => (x"71",x"7e",x"74",x"49"),
   320 => (x"87",x"cd",x"05",x"99"),
   321 => (x"c1",x"49",x"66",x"cc"),
   322 => (x"71",x"7e",x"74",x"99"),
   323 => (x"c4",x"c1",x"02",x"99"),
   324 => (x"4c",x"c8",x"ff",x"87"),
   325 => (x"cc",x"4b",x"66",x"c8"),
   326 => (x"bf",x"ec",x"48",x"a6"),
   327 => (x"87",x"fa",x"e2",x"78"),
   328 => (x"6c",x"5b",x"a6",x"cc"),
   329 => (x"d4",x"88",x"73",x"48"),
   330 => (x"e8",x"cf",x"58",x"a6"),
   331 => (x"87",x"d1",x"06",x"a8"),
   332 => (x"bf",x"fc",x"de",x"c2"),
   333 => (x"c2",x"b9",x"c1",x"49"),
   334 => (x"71",x"59",x"c0",x"df"),
   335 => (x"6c",x"87",x"c9",x"fd"),
   336 => (x"e7",x"49",x"c7",x"4b"),
   337 => (x"98",x"70",x"87",x"d1"),
   338 => (x"87",x"cb",x"ff",x"05"),
   339 => (x"c1",x"49",x"66",x"cc"),
   340 => (x"c2",x"ff",x"05",x"99"),
   341 => (x"c2",x"4c",x"6e",x"87"),
   342 => (x"4a",x"bf",x"c8",x"df"),
   343 => (x"df",x"c2",x"ba",x"c1"),
   344 => (x"0a",x"fc",x"5a",x"cc"),
   345 => (x"9a",x"c1",x"0a",x"7a"),
   346 => (x"49",x"a2",x"c0",x"c1"),
   347 => (x"c1",x"87",x"c7",x"e9"),
   348 => (x"e2",x"e6",x"49",x"da"),
   349 => (x"48",x"a6",x"c8",x"87"),
   350 => (x"df",x"c2",x"78",x"c1"),
   351 => (x"66",x"cc",x"48",x"c0"),
   352 => (x"c8",x"df",x"c2",x"78"),
   353 => (x"c7",x"c1",x"05",x"bf"),
   354 => (x"c0",x"c0",x"c8",x"87"),
   355 => (x"ec",x"de",x"c2",x"4b"),
   356 => (x"14",x"4c",x"6e",x"7e"),
   357 => (x"87",x"ff",x"e5",x"49"),
   358 => (x"c0",x"02",x"98",x"70"),
   359 => (x"b5",x"73",x"87",x"c2"),
   360 => (x"05",x"2b",x"b7",x"c1"),
   361 => (x"75",x"87",x"ec",x"ff"),
   362 => (x"99",x"ff",x"c3",x"49"),
   363 => (x"49",x"c0",x"1e",x"71"),
   364 => (x"75",x"87",x"c6",x"fb"),
   365 => (x"29",x"b7",x"c8",x"49"),
   366 => (x"49",x"c1",x"1e",x"71"),
   367 => (x"c8",x"87",x"fa",x"fa"),
   368 => (x"49",x"fd",x"c3",x"86"),
   369 => (x"c3",x"87",x"d0",x"e5"),
   370 => (x"ca",x"e5",x"49",x"fa"),
   371 => (x"87",x"ce",x"c7",x"87"),
   372 => (x"ff",x"c3",x"49",x"75"),
   373 => (x"2d",x"b7",x"c8",x"99"),
   374 => (x"9d",x"75",x"b5",x"71"),
   375 => (x"87",x"e0",x"c0",x"02"),
   376 => (x"7e",x"bf",x"c8",x"ff"),
   377 => (x"df",x"c2",x"49",x"6e"),
   378 => (x"c2",x"89",x"bf",x"c4"),
   379 => (x"c0",x"03",x"a9",x"e0"),
   380 => (x"4d",x"c0",x"87",x"c5"),
   381 => (x"c2",x"87",x"cf",x"c0"),
   382 => (x"6e",x"48",x"c4",x"df"),
   383 => (x"87",x"c6",x"c0",x"78"),
   384 => (x"48",x"c4",x"df",x"c2"),
   385 => (x"49",x"75",x"78",x"c0"),
   386 => (x"c0",x"05",x"99",x"c8"),
   387 => (x"f5",x"c3",x"87",x"ce"),
   388 => (x"87",x"c3",x"e4",x"49"),
   389 => (x"99",x"c2",x"49",x"70"),
   390 => (x"87",x"ea",x"c0",x"02"),
   391 => (x"bf",x"cc",x"fb",x"c2"),
   392 => (x"87",x"ca",x"c0",x"02"),
   393 => (x"c2",x"88",x"c1",x"48"),
   394 => (x"c0",x"58",x"d0",x"fb"),
   395 => (x"66",x"c4",x"87",x"d3"),
   396 => (x"80",x"e0",x"c1",x"48"),
   397 => (x"bf",x"6e",x"7e",x"70"),
   398 => (x"87",x"c5",x"c0",x"02"),
   399 => (x"73",x"49",x"ff",x"4b"),
   400 => (x"48",x"a6",x"c8",x"0f"),
   401 => (x"49",x"75",x"78",x"c1"),
   402 => (x"c0",x"05",x"99",x"c4"),
   403 => (x"f2",x"c3",x"87",x"ce"),
   404 => (x"87",x"c3",x"e3",x"49"),
   405 => (x"99",x"c2",x"49",x"70"),
   406 => (x"87",x"f1",x"c0",x"02"),
   407 => (x"bf",x"cc",x"fb",x"c2"),
   408 => (x"c7",x"48",x"6e",x"7e"),
   409 => (x"c0",x"03",x"a8",x"b7"),
   410 => (x"48",x"6e",x"87",x"cb"),
   411 => (x"fb",x"c2",x"80",x"c1"),
   412 => (x"d3",x"c0",x"58",x"d0"),
   413 => (x"48",x"66",x"c4",x"87"),
   414 => (x"70",x"80",x"e0",x"c1"),
   415 => (x"02",x"bf",x"6e",x"7e"),
   416 => (x"4b",x"87",x"c5",x"c0"),
   417 => (x"0f",x"73",x"49",x"fe"),
   418 => (x"c1",x"48",x"a6",x"c8"),
   419 => (x"49",x"fd",x"c3",x"78"),
   420 => (x"70",x"87",x"c4",x"e2"),
   421 => (x"02",x"99",x"c2",x"49"),
   422 => (x"c2",x"87",x"e6",x"c0"),
   423 => (x"02",x"bf",x"cc",x"fb"),
   424 => (x"c2",x"87",x"c9",x"c0"),
   425 => (x"c0",x"48",x"cc",x"fb"),
   426 => (x"87",x"d0",x"c0",x"78"),
   427 => (x"c1",x"4a",x"66",x"c4"),
   428 => (x"02",x"6a",x"82",x"e0"),
   429 => (x"4b",x"87",x"c5",x"c0"),
   430 => (x"0f",x"73",x"49",x"fd"),
   431 => (x"c1",x"48",x"a6",x"c8"),
   432 => (x"49",x"fa",x"c3",x"78"),
   433 => (x"70",x"87",x"d0",x"e1"),
   434 => (x"02",x"99",x"c2",x"49"),
   435 => (x"c2",x"87",x"ed",x"c0"),
   436 => (x"48",x"bf",x"cc",x"fb"),
   437 => (x"03",x"a8",x"b7",x"c7"),
   438 => (x"c2",x"87",x"c9",x"c0"),
   439 => (x"c7",x"48",x"cc",x"fb"),
   440 => (x"87",x"d3",x"c0",x"78"),
   441 => (x"c1",x"48",x"66",x"c4"),
   442 => (x"7e",x"70",x"80",x"e0"),
   443 => (x"c0",x"02",x"bf",x"6e"),
   444 => (x"fc",x"4b",x"87",x"c5"),
   445 => (x"c8",x"0f",x"73",x"49"),
   446 => (x"78",x"c1",x"48",x"a6"),
   447 => (x"f0",x"c3",x"48",x"75"),
   448 => (x"48",x"7e",x"70",x"98"),
   449 => (x"ce",x"c0",x"05",x"98"),
   450 => (x"49",x"da",x"c1",x"87"),
   451 => (x"70",x"87",x"c8",x"e0"),
   452 => (x"02",x"99",x"c2",x"49"),
   453 => (x"6e",x"87",x"ca",x"c1"),
   454 => (x"87",x"cd",x"c0",x"05"),
   455 => (x"ff",x"49",x"da",x"c1"),
   456 => (x"70",x"87",x"f4",x"df"),
   457 => (x"e8",x"c0",x"02",x"98"),
   458 => (x"49",x"bf",x"e8",x"87"),
   459 => (x"9b",x"ff",x"c3",x"4b"),
   460 => (x"71",x"29",x"b7",x"c8"),
   461 => (x"e1",x"da",x"ff",x"b3"),
   462 => (x"c3",x"49",x"73",x"87"),
   463 => (x"99",x"71",x"99",x"f0"),
   464 => (x"87",x"e5",x"ff",x"05"),
   465 => (x"ff",x"49",x"da",x"c1"),
   466 => (x"70",x"87",x"cc",x"df"),
   467 => (x"d8",x"ff",x"05",x"98"),
   468 => (x"cc",x"fb",x"c2",x"87"),
   469 => (x"cc",x"4b",x"49",x"bf"),
   470 => (x"83",x"66",x"c4",x"93"),
   471 => (x"73",x"71",x"4b",x"6b"),
   472 => (x"02",x"9c",x"74",x"0f"),
   473 => (x"6c",x"87",x"e9",x"c0"),
   474 => (x"87",x"e4",x"c0",x"02"),
   475 => (x"de",x"ff",x"49",x"6c"),
   476 => (x"49",x"70",x"87",x"e5"),
   477 => (x"c0",x"02",x"99",x"c1"),
   478 => (x"a4",x"c4",x"87",x"cb"),
   479 => (x"cc",x"fb",x"c2",x"4b"),
   480 => (x"4b",x"6b",x"49",x"bf"),
   481 => (x"02",x"84",x"c8",x"0f"),
   482 => (x"6c",x"87",x"c5",x"c0"),
   483 => (x"87",x"dc",x"ff",x"05"),
   484 => (x"c0",x"02",x"66",x"c8"),
   485 => (x"fb",x"c2",x"87",x"c8"),
   486 => (x"f1",x"49",x"bf",x"cc"),
   487 => (x"8e",x"ec",x"87",x"de"),
   488 => (x"4c",x"26",x"4d",x"26"),
   489 => (x"4f",x"26",x"4b",x"26"),
   490 => (x"00",x"00",x"00",x"10"),
   491 => (x"14",x"11",x"12",x"58"),
   492 => (x"23",x"1c",x"1b",x"1d"),
   493 => (x"94",x"91",x"59",x"5a"),
   494 => (x"f4",x"eb",x"f2",x"f5"),
   495 => (x"00",x"00",x"00",x"00"),
   496 => (x"00",x"00",x"00",x"00"),
   497 => (x"00",x"00",x"00",x"00"),
   498 => (x"00",x"00",x"00",x"00"),
   499 => (x"5c",x"5b",x"5e",x"0e"),
   500 => (x"4b",x"71",x"0e",x"5d"),
   501 => (x"d0",x"4c",x"d4",x"ff"),
   502 => (x"78",x"c0",x"48",x"66"),
   503 => (x"dd",x"ff",x"49",x"d6"),
   504 => (x"ff",x"c3",x"87",x"f2"),
   505 => (x"c3",x"49",x"6c",x"7c"),
   506 => (x"4d",x"71",x"99",x"ff"),
   507 => (x"99",x"f0",x"c3",x"49"),
   508 => (x"05",x"a9",x"e0",x"c1"),
   509 => (x"ff",x"c3",x"87",x"cb"),
   510 => (x"c3",x"48",x"6c",x"7c"),
   511 => (x"08",x"66",x"d0",x"98"),
   512 => (x"7c",x"ff",x"c3",x"78"),
   513 => (x"c8",x"49",x"4a",x"6c"),
   514 => (x"7c",x"ff",x"c3",x"31"),
   515 => (x"b2",x"71",x"4a",x"6c"),
   516 => (x"31",x"c8",x"49",x"72"),
   517 => (x"6c",x"7c",x"ff",x"c3"),
   518 => (x"72",x"b2",x"71",x"4a"),
   519 => (x"c3",x"31",x"c8",x"49"),
   520 => (x"4a",x"6c",x"7c",x"ff"),
   521 => (x"d0",x"ff",x"b2",x"71"),
   522 => (x"78",x"e0",x"c0",x"48"),
   523 => (x"c2",x"02",x"9b",x"73"),
   524 => (x"75",x"7b",x"72",x"87"),
   525 => (x"26",x"4d",x"26",x"48"),
   526 => (x"26",x"4b",x"26",x"4c"),
   527 => (x"4f",x"26",x"1e",x"4f"),
   528 => (x"5c",x"5b",x"5e",x"0e"),
   529 => (x"76",x"86",x"f8",x"0e"),
   530 => (x"49",x"a6",x"c8",x"1e"),
   531 => (x"c4",x"87",x"fd",x"fd"),
   532 => (x"6e",x"4b",x"70",x"86"),
   533 => (x"01",x"a8",x"c3",x"48"),
   534 => (x"73",x"87",x"f4",x"c2"),
   535 => (x"9a",x"f0",x"c3",x"4a"),
   536 => (x"02",x"aa",x"d0",x"c1"),
   537 => (x"e0",x"c1",x"87",x"c7"),
   538 => (x"e2",x"c2",x"05",x"aa"),
   539 => (x"c8",x"49",x"73",x"87"),
   540 => (x"87",x"c3",x"02",x"99"),
   541 => (x"73",x"87",x"c6",x"ff"),
   542 => (x"c2",x"9c",x"c3",x"4c"),
   543 => (x"c4",x"c1",x"05",x"ac"),
   544 => (x"49",x"66",x"c4",x"87"),
   545 => (x"1e",x"71",x"31",x"c9"),
   546 => (x"c1",x"4a",x"66",x"c4"),
   547 => (x"fb",x"c2",x"92",x"cc"),
   548 => (x"81",x"72",x"49",x"d4"),
   549 => (x"87",x"d6",x"cd",x"fe"),
   550 => (x"da",x"ff",x"49",x"d8"),
   551 => (x"c0",x"c8",x"87",x"f6"),
   552 => (x"cc",x"e8",x"c2",x"1e"),
   553 => (x"ec",x"e6",x"fd",x"49"),
   554 => (x"48",x"d0",x"ff",x"87"),
   555 => (x"c2",x"78",x"e0",x"c0"),
   556 => (x"cc",x"1e",x"cc",x"e8"),
   557 => (x"cc",x"c1",x"4a",x"66"),
   558 => (x"d4",x"fb",x"c2",x"92"),
   559 => (x"fe",x"81",x"72",x"49"),
   560 => (x"cc",x"87",x"ec",x"cb"),
   561 => (x"05",x"ac",x"c1",x"86"),
   562 => (x"c4",x"87",x"c4",x"c1"),
   563 => (x"31",x"c9",x"49",x"66"),
   564 => (x"66",x"c4",x"1e",x"71"),
   565 => (x"92",x"cc",x"c1",x"4a"),
   566 => (x"49",x"d4",x"fb",x"c2"),
   567 => (x"cc",x"fe",x"81",x"72"),
   568 => (x"e8",x"c2",x"87",x"cc"),
   569 => (x"66",x"c8",x"1e",x"cc"),
   570 => (x"92",x"cc",x"c1",x"4a"),
   571 => (x"49",x"d4",x"fb",x"c2"),
   572 => (x"c9",x"fe",x"81",x"72"),
   573 => (x"49",x"d7",x"87",x"fa"),
   574 => (x"87",x"d8",x"d9",x"ff"),
   575 => (x"c2",x"1e",x"c0",x"c8"),
   576 => (x"fd",x"49",x"cc",x"e8"),
   577 => (x"cc",x"87",x"eb",x"e4"),
   578 => (x"48",x"d0",x"ff",x"86"),
   579 => (x"f8",x"78",x"e0",x"c0"),
   580 => (x"26",x"4c",x"26",x"8e"),
   581 => (x"1e",x"4f",x"26",x"4b"),
   582 => (x"b7",x"c4",x"4a",x"71"),
   583 => (x"87",x"ce",x"03",x"aa"),
   584 => (x"cc",x"c1",x"49",x"72"),
   585 => (x"d4",x"fb",x"c2",x"91"),
   586 => (x"81",x"c8",x"c1",x"81"),
   587 => (x"4f",x"26",x"79",x"c0"),
   588 => (x"5c",x"5b",x"5e",x"0e"),
   589 => (x"86",x"fc",x"0e",x"5d"),
   590 => (x"d4",x"ff",x"4a",x"71"),
   591 => (x"d4",x"4c",x"c0",x"4b"),
   592 => (x"b7",x"c3",x"4d",x"66"),
   593 => (x"c2",x"c2",x"01",x"ad"),
   594 => (x"02",x"9a",x"72",x"87"),
   595 => (x"1e",x"87",x"ec",x"c0"),
   596 => (x"cc",x"c1",x"49",x"75"),
   597 => (x"d4",x"fb",x"c2",x"91"),
   598 => (x"c8",x"80",x"71",x"48"),
   599 => (x"66",x"c4",x"58",x"a6"),
   600 => (x"d7",x"c3",x"fe",x"49"),
   601 => (x"70",x"86",x"c4",x"87"),
   602 => (x"87",x"d4",x"02",x"98"),
   603 => (x"c8",x"c1",x"49",x"6e"),
   604 => (x"6e",x"79",x"c1",x"81"),
   605 => (x"69",x"81",x"c8",x"49"),
   606 => (x"75",x"87",x"c5",x"4c"),
   607 => (x"87",x"d7",x"fe",x"49"),
   608 => (x"c8",x"48",x"d0",x"ff"),
   609 => (x"7b",x"dd",x"78",x"e1"),
   610 => (x"ff",x"c3",x"48",x"74"),
   611 => (x"74",x"7b",x"70",x"98"),
   612 => (x"29",x"b7",x"c8",x"49"),
   613 => (x"ff",x"c3",x"48",x"71"),
   614 => (x"74",x"7b",x"70",x"98"),
   615 => (x"29",x"b7",x"d0",x"49"),
   616 => (x"ff",x"c3",x"48",x"71"),
   617 => (x"74",x"7b",x"70",x"98"),
   618 => (x"28",x"b7",x"d8",x"48"),
   619 => (x"7b",x"c0",x"7b",x"70"),
   620 => (x"7b",x"7b",x"7b",x"7b"),
   621 => (x"7b",x"7b",x"7b",x"7b"),
   622 => (x"ff",x"7b",x"7b",x"7b"),
   623 => (x"e0",x"c0",x"48",x"d0"),
   624 => (x"dc",x"1e",x"75",x"78"),
   625 => (x"f0",x"d6",x"ff",x"49"),
   626 => (x"fc",x"86",x"c4",x"87"),
   627 => (x"26",x"4d",x"26",x"8e"),
   628 => (x"26",x"4b",x"26",x"4c"),
   629 => (x"00",x"1c",x"ff",x"4f"),
   630 => (x"00",x"1c",x"ff",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

